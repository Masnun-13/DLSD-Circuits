CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 0 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
144
13 Logic Switch~
5 38 474 0 10 11
0 73 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
1 F
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44105.3 0
0
13 Logic Switch~
5 40 411 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
1 E
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44105.3 1
0
13 Logic Switch~
5 43 369 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -17 8 -9
1 D
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
44105.3 2
0
13 Logic Switch~
5 67 163 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-9 -15 5 -7
1 C
-4 -29 3 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44105.3 3
0
13 Logic Switch~
5 66 214 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44105.3 4
0
13 Logic Switch~
5 63 263 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -17 8 -9
1 A
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
44105.3 5
0
9 Inverter~
13 1639 543 0 2 22
0 9 10
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
8901 0 0
2
44105.3 6
0
14 Logic Display~
6 1642 509 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out63
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
44105.3 7
0
9 Inverter~
13 1592 542 0 2 22
0 11 12
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
4747 0 0
2
44105.3 8
0
14 Logic Display~
6 1595 508 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out62
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
44105.3 9
0
9 Inverter~
13 1547 543 0 2 22
0 13 14
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 6 0
1 U
3472 0 0
2
44105.3 10
0
14 Logic Display~
6 1550 509 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out61
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
44105.3 11
0
9 Inverter~
13 1497 545 0 2 22
0 15 16
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
3536 0 0
2
44105.3 12
0
14 Logic Display~
6 1500 511 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out60
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44105.3 13
0
9 Inverter~
13 1443 542 0 2 22
0 17 18
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
3835 0 0
2
44105.3 14
0
14 Logic Display~
6 1446 508 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out59
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
44105.3 15
0
9 Inverter~
13 1397 543 0 2 22
0 19 20
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
5616 0 0
2
44105.3 16
0
14 Logic Display~
6 1400 509 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out58
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
44105.3 17
0
9 Inverter~
13 1348 542 0 2 22
0 21 22
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 7 0
1 U
317 0 0
2
44105.3 18
0
14 Logic Display~
6 1351 508 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out57
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44105.3 19
0
9 Inverter~
13 1305 540 0 2 22
0 23 24
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 7 0
1 U
4299 0 0
2
44105.3 20
0
14 Logic Display~
6 1308 506 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out56
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
44105.3 21
0
9 Inverter~
13 1639 406 0 2 22
0 25 26
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 7 0
1 U
7876 0 0
2
44105.3 22
0
14 Logic Display~
6 1642 372 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out55
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
44105.3 23
0
9 Inverter~
13 1592 405 0 2 22
0 27 28
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
9172 0 0
2
44105.3 24
0
14 Logic Display~
6 1595 371 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out54
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
44105.3 25
0
9 Inverter~
13 1549 404 0 2 22
0 29 30
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
3820 0 0
2
44105.3 26
0
14 Logic Display~
6 1552 370 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out53
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
44105.3 27
0
9 Inverter~
13 1498 406 0 2 22
0 31 32
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
961 0 0
2
44105.3 28
0
14 Logic Display~
6 1501 372 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out52
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
44105.3 29
0
9 Inverter~
13 1444 407 0 2 22
0 33 34
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
3409 0 0
2
44105.3 30
0
14 Logic Display~
6 1447 373 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out51
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
44105.3 31
0
9 Inverter~
13 1398 406 0 2 22
0 35 36
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
8885 0 0
2
44105.3 32
0
14 Logic Display~
6 1401 372 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out50
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
44105.3 33
0
9 Inverter~
13 1349 406 0 2 22
0 37 38
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
9265 0 0
2
44105.3 34
0
14 Logic Display~
6 1352 372 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out49
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
44105.3 35
0
9 Inverter~
13 1306 407 0 2 22
0 39 40
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
9424 0 0
2
44105.3 36
0
14 Logic Display~
6 1309 373 0 1 2
10 40
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out48
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
44105.3 37
0
9 Inverter~
13 1635 270 0 2 22
0 41 42
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
9281 0 0
2
44105.3 38
0
14 Logic Display~
6 1638 236 0 1 2
10 42
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out47
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
44105.3 39
0
9 Inverter~
13 1588 268 0 2 22
0 43 44
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
7168 0 0
2
44105.3 40
0
14 Logic Display~
6 1591 234 0 1 2
10 44
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out46
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
44105.3 41
0
9 Inverter~
13 1545 268 0 2 22
0 45 46
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
4139 0 0
2
44105.3 42
0
14 Logic Display~
6 1548 234 0 1 2
10 46
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out45
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
44105.3 43
0
9 Inverter~
13 1494 269 0 2 22
0 47 48
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
5283 0 0
2
44105.3 44
0
14 Logic Display~
6 1497 235 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out44
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
44105.3 45
0
9 Inverter~
13 1440 267 0 2 22
0 49 50
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
5305 0 0
2
44105.3 46
0
14 Logic Display~
6 1443 233 0 1 2
10 50
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out43
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
44105.3 47
0
9 Inverter~
13 1394 267 0 2 22
0 51 52
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
969 0 0
2
44105.3 48
0
14 Logic Display~
6 1397 233 0 1 2
10 52
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out42
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
44105.3 49
0
9 Inverter~
13 1345 267 0 2 22
0 53 54
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
3751 0 0
2
44105.3 50
0
14 Logic Display~
6 1348 233 0 1 2
10 54
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out41
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
44105.3 51
0
9 Inverter~
13 1300 265 0 2 22
0 55 56
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
6118 0 0
2
44105.3 52
0
14 Logic Display~
6 1303 231 0 1 2
10 56
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out40
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
44105.3 53
0
9 Inverter~
13 1636 123 0 2 22
0 57 58
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
6357 0 0
2
44105.3 54
0
14 Logic Display~
6 1639 89 0 1 2
10 58
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out39
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
44105.3 55
0
9 Inverter~
13 1589 115 0 2 22
0 70 59
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
3976 0 0
2
44105.3 56
0
14 Logic Display~
6 1592 81 0 1 2
10 59
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out38
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
44105.3 57
0
9 Inverter~
13 1546 118 0 2 22
0 60 61
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
523 0 0
2
44105.3 58
0
14 Logic Display~
6 1549 84 0 1 2
10 61
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out37
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
44105.3 59
0
9 Inverter~
13 1495 120 0 2 22
0 62 63
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
6901 0 0
2
44105.3 60
0
14 Logic Display~
6 1498 86 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out36
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
44105.3 61
0
9 Inverter~
13 1441 119 0 2 22
0 64 65
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
3277 0 0
2
44105.3 62
0
14 Logic Display~
6 1444 85 0 1 2
10 65
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Ou35
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
44105.3 63
0
9 Inverter~
13 1395 118 0 2 22
0 71 66
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
4720 0 0
2
44105.3 64
0
14 Logic Display~
6 1398 84 0 1 2
10 66
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out34
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5551 0 0
2
44105.3 65
0
9 Inverter~
13 1346 120 0 2 22
0 72 67
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
6986 0 0
2
44105.3 66
0
14 Logic Display~
6 1349 86 0 1 2
10 67
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out33
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8745 0 0
2
44105.3 67
0
14 Logic Display~
6 1303 86 0 1 2
10 68
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out32
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
44105.3 68
0
9 Inverter~
13 1300 120 0 2 22
0 69 68
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 11 0
1 U
8748 0 0
2
44105.3 69
0
7 74LS138
19 1224 184 0 14 29
0 7 6 5 8 3 2 57 70 60
62 64 71 72 69
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U16
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7168 0 0
2
44105.3 70
0
7 74LS138
19 1233 597 0 14 29
0 7 6 5 3 8 2 9 11 13
15 17 19 21 23
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U17
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
631 0 0
2
44105.3 71
0
7 74LS138
19 1229 459 0 14 29
0 7 6 5 3 4 2 25 27 29
31 33 35 37 39
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U18
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
9466 0 0
2
44105.3 72
0
7 74LS138
19 1228 328 0 14 29
0 7 6 5 4 3 2 41 43 45
47 49 51 53 55
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U19
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3266 0 0
2
44105.3 73
0
9 Inverter~
13 886 529 0 2 22
0 73 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 11 0
1 U
7693 0 0
2
44105.3 74
0
9 Inverter~
13 740 549 0 2 22
0 74 75
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
3723 0 0
2
44105.3 75
0
14 Logic Display~
6 743 515 0 1 2
10 75
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out31
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
44105.3 76
0
9 Inverter~
13 693 548 0 2 22
0 76 77
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
6263 0 0
2
44105.3 77
0
14 Logic Display~
6 696 514 0 1 2
10 77
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out30
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4900 0 0
2
44105.3 78
0
9 Inverter~
13 648 549 0 2 22
0 78 79
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
8783 0 0
2
44105.3 79
0
14 Logic Display~
6 651 515 0 1 2
10 79
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out29
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3221 0 0
2
44105.3 80
0
9 Inverter~
13 598 551 0 2 22
0 80 81
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 5 0
1 U
3215 0 0
2
44105.3 81
0
14 Logic Display~
6 601 517 0 1 2
10 81
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out28
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
44105.3 82
0
9 Inverter~
13 544 548 0 2 22
0 82 83
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 5 0
1 U
7121 0 0
2
44105.3 83
0
14 Logic Display~
6 547 514 0 1 2
10 83
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out27
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
44105.3 84
0
9 Inverter~
13 498 549 0 2 22
0 84 85
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
5996 0 0
2
44105.3 85
0
14 Logic Display~
6 501 515 0 1 2
10 85
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out26
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7804 0 0
2
44105.3 86
0
9 Inverter~
13 449 548 0 2 22
0 86 87
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
5523 0 0
2
44105.3 87
0
14 Logic Display~
6 452 514 0 1 2
10 87
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out25
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
44105.3 88
0
9 Inverter~
13 406 546 0 2 22
0 88 89
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
3465 0 0
2
44105.3 89
0
14 Logic Display~
6 409 512 0 1 2
10 89
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out24
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
44105.3 90
0
9 Inverter~
13 740 412 0 2 22
0 90 91
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3685 0 0
2
44105.3 91
0
14 Logic Display~
6 743 378 0 1 2
10 91
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out23
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
44105.3 92
0
9 Inverter~
13 693 411 0 2 22
0 92 93
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
6343 0 0
2
44105.3 93
0
14 Logic Display~
6 696 377 0 1 2
10 93
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out22
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
44105.3 94
0
9 Inverter~
13 650 410 0 2 22
0 94 95
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
9156 0 0
2
44105.3 95
0
14 Logic Display~
6 653 376 0 1 2
10 95
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out21
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
44105.3 96
0
9 Inverter~
13 599 412 0 2 22
0 96 97
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
7207 0 0
2
44105.3 97
0
14 Logic Display~
6 602 378 0 1 2
10 97
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out20
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
44105.3 98
0
9 Inverter~
13 545 413 0 2 22
0 98 99
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
3760 0 0
2
44105.3 99
0
14 Logic Display~
6 548 379 0 1 2
10 99
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out19
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
44105.3 100
0
9 Inverter~
13 499 412 0 2 22
0 100 101
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9767 0 0
2
44105.3 101
0
14 Logic Display~
6 502 378 0 1 2
10 101
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out18
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7978 0 0
2
44105.3 102
0
9 Inverter~
13 450 412 0 2 22
0 102 103
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3142 0 0
2
44105.3 103
0
14 Logic Display~
6 453 378 0 1 2
10 103
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out17
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3284 0 0
2
44105.3 104
0
9 Inverter~
13 407 413 0 2 22
0 104 105
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
659 0 0
2
44105.3 105
0
14 Logic Display~
6 410 379 0 1 2
10 105
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out16
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
44105.3 106
0
9 Inverter~
13 736 276 0 2 22
0 106 107
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
6792 0 0
2
44105.3 107
0
14 Logic Display~
6 739 242 0 1 2
10 107
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out15
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
44105.3 108
0
9 Inverter~
13 689 274 0 2 22
0 108 109
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
6316 0 0
2
44105.3 109
0
14 Logic Display~
6 692 240 0 1 2
10 109
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out14
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8734 0 0
2
44105.3 110
0
9 Inverter~
13 646 274 0 2 22
0 110 111
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
7988 0 0
2
44105.3 111
0
14 Logic Display~
6 649 240 0 1 2
10 111
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out13
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3217 0 0
2
44105.3 112
0
9 Inverter~
13 595 275 0 2 22
0 112 113
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3965 0 0
2
44105.3 113
0
14 Logic Display~
6 598 241 0 1 2
10 113
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out12
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8239 0 0
2
44105.3 114
0
9 Inverter~
13 541 273 0 2 22
0 114 115
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
828 0 0
2
44105.3 115
0
14 Logic Display~
6 544 239 0 1 2
10 115
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out11
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
44105.3 116
0
9 Inverter~
13 495 273 0 2 22
0 116 117
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
7107 0 0
2
44105.3 117
0
14 Logic Display~
6 498 239 0 1 2
10 117
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out10
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6433 0 0
2
44105.3 118
0
9 Inverter~
13 446 273 0 2 22
0 118 119
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
8559 0 0
2
44105.3 119
0
14 Logic Display~
6 449 239 0 1 2
10 119
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out9
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3674 0 0
2
44105.3 120
0
9 Inverter~
13 401 271 0 2 22
0 120 121
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
5697 0 0
2
44105.3 121
0
14 Logic Display~
6 404 237 0 1 2
10 121
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out8
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3805 0 0
2
44105.3 122
0
9 Inverter~
13 737 129 0 2 22
0 122 123
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
5219 0 0
2
44105.3 123
0
14 Logic Display~
6 740 95 0 1 2
10 123
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out7
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3795 0 0
2
44105.3 124
0
9 Inverter~
13 690 121 0 2 22
0 135 124
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3637 0 0
2
44105.3 125
0
14 Logic Display~
6 693 87 0 1 2
10 124
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out6
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
44105.3 126
0
9 Inverter~
13 647 124 0 2 22
0 125 126
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6966 0 0
2
44105.3 127
0
14 Logic Display~
6 650 90 0 1 2
10 126
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out5
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9796 0 0
2
44105.3 128
0
9 Inverter~
13 596 126 0 2 22
0 127 128
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
5952 0 0
2
44105.3 129
0
14 Logic Display~
6 599 92 0 1 2
10 128
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out4
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3649 0 0
2
44105.3 130
0
9 Inverter~
13 542 125 0 2 22
0 129 130
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3716 0 0
2
44105.3 131
0
14 Logic Display~
6 545 91 0 1 2
10 130
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out3
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
44105.3 132
0
9 Inverter~
13 496 124 0 2 22
0 136 131
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4681 0 0
2
44105.3 133
0
14 Logic Display~
6 499 90 0 1 2
10 131
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out2
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9730 0 0
2
44105.3 134
0
9 Inverter~
13 447 126 0 2 22
0 137 132
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9874 0 0
2
44105.3 135
0
14 Logic Display~
6 450 92 0 1 2
10 132
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out1
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
364 0 0
2
44105.3 136
0
14 Logic Display~
6 404 92 0 1 2
10 133
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out00
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3656 0 0
2
44105.3 137
0
9 Inverter~
13 401 126 0 2 22
0 134 133
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3131 0 0
2
44105.3 138
0
9 Inverter~
13 77 346 0 2 22
0 4 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6772 0 0
2
44105.3 139
0
7 74LS138
19 332 189 0 14 29
0 7 6 5 8 73 3 122 135 125
127 129 136 137 134
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
9557 0 0
2
44105.3 140
0
7 74LS138
19 334 603 0 14 29
0 7 6 5 3 8 73 74 76 78
80 82 84 86 88
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U4
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
5789 0 0
2
44105.3 141
0
7 74LS138
19 330 465 0 14 29
0 7 6 5 3 4 73 90 92 94
96 98 100 102 104
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U3
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7328 0 0
2
44105.3 142
0
7 74LS138
19 331 335 0 14 29
0 7 6 5 4 3 73 106 108 110
112 114 116 118 120
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U2
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
4799 0 0
2
44105.3 143
0
258
6 0 2 0 0 4096 0 74 0 0 123 4
1190 364
1196 364
1196 364
1192 364
5 0 3 0 0 4096 0 74 0 0 120 4
1190 355
1196 355
1196 355
1192 355
4 0 4 0 0 4096 0 74 0 0 128 4
1196 346
1202 346
1202 346
1198 346
3 0 5 0 0 4096 0 74 0 0 132 4
1196 319
1202 319
1202 319
1198 319
2 0 6 0 0 4096 0 74 0 0 136 4
1196 310
1202 310
1202 310
1198 310
1 0 7 0 0 4096 0 74 0 0 140 4
1196 301
1202 301
1202 301
1198 301
6 0 2 0 0 0 0 73 0 0 124 2
1191 495
1191 494
5 0 4 0 0 0 0 73 0 0 119 2
1191 486
1191 485
4 0 3 0 0 0 0 73 0 0 127 2
1197 477
1197 476
3 0 5 0 0 0 0 73 0 0 131 2
1197 450
1197 449
2 0 6 0 0 0 0 73 0 0 135 2
1197 441
1197 440
1 0 7 0 0 0 0 73 0 0 139 2
1197 432
1197 431
6 0 2 0 0 0 0 72 0 0 125 2
1195 633
1195 632
5 0 8 0 0 4096 0 72 0 0 118 2
1195 624
1195 623
4 0 3 0 0 0 0 72 0 0 117 2
1201 615
1201 614
3 0 5 0 0 0 0 72 0 0 130 2
1201 588
1201 587
2 0 6 0 0 0 0 72 0 0 134 2
1201 579
1201 578
1 0 7 0 0 0 0 72 0 0 138 2
1201 570
1201 569
6 0 2 0 0 8192 0 71 0 0 122 3
1186 220
1186 218
1193 218
5 0 3 0 0 8192 0 71 0 0 121 3
1186 211
1186 209
1193 209
4 0 8 0 0 8192 0 71 0 0 129 3
1192 202
1192 200
1199 200
3 0 5 0 0 8192 0 71 0 0 133 3
1192 175
1192 173
1199 173
2 0 6 0 0 8192 0 71 0 0 137 3
1192 166
1192 164
1199 164
1 0 7 0 0 8192 0 71 0 0 141 3
1192 157
1192 155
1199 155
1 0 9 0 0 4096 0 7 0 0 94 2
1642 561
1641 561
1 2 10 0 0 4224 0 8 7 0 0 2
1642 527
1642 525
1 0 11 0 0 4096 0 9 0 0 95 2
1595 560
1594 560
1 2 12 0 0 4224 0 10 9 0 0 2
1595 526
1595 524
1 0 13 0 0 4096 0 11 0 0 86 2
1550 561
1551 561
1 2 14 0 0 4224 0 12 11 0 0 2
1550 527
1550 525
1 0 15 0 0 0 0 13 0 0 96 2
1500 563
1500 563
1 2 16 0 0 4224 0 14 13 0 0 2
1500 529
1500 527
1 0 17 0 0 0 0 15 0 0 97 2
1446 560
1446 560
1 2 18 0 0 4224 0 16 15 0 0 2
1446 526
1446 524
1 0 19 0 0 0 0 17 0 0 98 2
1400 561
1400 561
1 2 20 0 0 4224 0 18 17 0 0 2
1400 527
1400 525
1 0 21 0 0 0 0 19 0 0 99 2
1351 560
1351 560
1 2 22 0 0 4224 0 20 19 0 0 2
1351 526
1351 524
1 0 23 0 0 0 0 21 0 0 100 2
1308 558
1308 558
1 2 24 0 0 4224 0 22 21 0 0 2
1308 524
1308 522
1 0 25 0 0 0 0 23 0 0 101 2
1642 424
1642 424
1 2 26 0 0 4224 0 24 23 0 0 2
1642 390
1642 388
1 0 27 0 0 0 0 25 0 0 102 2
1595 423
1595 423
1 2 28 0 0 4224 0 26 25 0 0 2
1595 389
1595 387
1 0 29 0 0 0 0 27 0 0 103 2
1552 422
1552 422
1 2 30 0 0 4224 0 28 27 0 0 2
1552 388
1552 386
1 0 31 0 0 0 0 29 0 0 104 2
1501 424
1501 424
1 2 32 0 0 4224 0 30 29 0 0 2
1501 390
1501 388
1 0 33 0 0 0 0 31 0 0 105 2
1447 425
1447 425
1 2 34 0 0 4224 0 32 31 0 0 2
1447 391
1447 389
1 0 35 0 0 0 0 33 0 0 106 2
1401 424
1401 424
1 2 36 0 0 4224 0 34 33 0 0 2
1401 390
1401 388
1 0 37 0 0 0 0 35 0 0 107 2
1352 424
1352 424
1 2 38 0 0 4224 0 36 35 0 0 2
1352 390
1352 388
1 0 39 0 0 0 0 37 0 0 108 2
1309 425
1309 425
1 2 40 0 0 4224 0 38 37 0 0 2
1309 391
1309 389
1 0 41 0 0 0 0 39 0 0 109 2
1638 288
1638 288
1 2 42 0 0 4224 0 40 39 0 0 2
1638 254
1638 252
1 0 43 0 0 0 0 41 0 0 110 2
1591 286
1591 286
1 2 44 0 0 4224 0 42 41 0 0 2
1591 252
1591 250
1 0 45 0 0 0 0 43 0 0 111 2
1548 286
1548 286
1 2 46 0 0 4224 0 44 43 0 0 2
1548 252
1548 250
1 0 47 0 0 0 0 45 0 0 112 2
1497 287
1497 287
1 2 48 0 0 4224 0 46 45 0 0 2
1497 253
1497 251
1 0 49 0 0 0 0 47 0 0 113 2
1443 285
1443 285
1 2 50 0 0 4224 0 48 47 0 0 2
1443 251
1443 249
1 0 51 0 0 0 0 49 0 0 114 2
1397 285
1397 285
1 2 52 0 0 4224 0 50 49 0 0 2
1397 251
1397 249
1 0 53 0 0 0 0 51 0 0 115 2
1348 285
1348 285
1 2 54 0 0 4224 0 52 51 0 0 2
1348 251
1348 249
1 0 55 0 0 0 0 53 0 0 116 2
1303 283
1303 283
1 2 56 0 0 4224 0 54 53 0 0 2
1303 249
1303 247
1 0 57 0 0 0 0 55 0 0 87 2
1639 141
1639 141
1 2 58 0 0 4224 0 56 55 0 0 2
1639 107
1639 105
1 2 59 0 0 4224 0 58 57 0 0 2
1592 99
1592 97
1 0 60 0 0 0 0 59 0 0 89 2
1549 136
1549 136
1 2 61 0 0 4224 0 60 59 0 0 2
1549 102
1549 100
1 0 62 0 0 0 0 61 0 0 90 2
1498 138
1498 138
1 2 63 0 0 4224 0 62 61 0 0 2
1498 104
1498 102
1 0 64 0 0 0 0 63 0 0 91 2
1444 137
1444 137
1 2 65 0 0 4224 0 64 63 0 0 2
1444 103
1444 101
1 2 66 0 0 4224 0 66 65 0 0 2
1398 102
1398 100
1 2 67 0 0 4224 0 68 67 0 0 2
1349 104
1349 102
1 2 68 0 0 4224 0 69 70 0 0 2
1303 104
1303 102
14 1 69 0 0 8320 0 71 70 0 0 3
1262 220
1303 220
1303 138
0 9 13 0 0 8320 0 0 72 0 0 3
1551 548
1551 588
1271 588
7 0 57 0 0 4224 0 71 0 0 0 3
1262 157
1639 157
1639 137
1 8 70 0 0 8320 0 57 71 0 0 3
1592 133
1592 166
1262 166
9 0 60 0 0 4224 0 71 0 0 0 3
1262 175
1549 175
1549 132
10 0 62 0 0 4224 0 71 0 0 0 3
1262 184
1498 184
1498 134
11 0 64 0 0 4224 0 71 0 0 0 3
1262 193
1444 193
1444 134
12 1 71 0 0 4224 0 71 65 0 0 3
1262 202
1398 202
1398 136
13 1 72 0 0 4224 0 71 67 0 0 3
1262 211
1349 211
1349 138
7 0 9 0 0 4224 0 72 0 0 0 3
1271 570
1641 570
1641 551
0 8 11 0 0 8320 0 0 72 0 0 3
1594 546
1594 579
1271 579
10 0 15 0 0 4224 0 72 0 0 0 3
1271 597
1500 597
1500 548
11 0 17 0 0 4224 0 72 0 0 0 3
1271 606
1446 606
1446 548
12 0 19 0 0 4224 0 72 0 0 0 3
1271 615
1400 615
1400 548
13 0 21 0 0 4224 0 72 0 0 0 3
1271 624
1351 624
1351 550
0 14 23 0 0 4224 0 0 72 0 0 3
1308 549
1308 633
1271 633
7 0 25 0 0 4224 0 73 0 0 0 3
1267 432
1642 432
1642 419
0 8 27 0 0 8320 0 0 73 0 0 3
1595 414
1595 441
1267 441
9 0 29 0 0 4224 0 73 0 0 0 3
1267 450
1552 450
1552 414
10 0 31 0 0 4224 0 73 0 0 0 3
1267 459
1501 459
1501 416
11 0 33 0 0 4224 0 73 0 0 0 3
1267 468
1447 468
1447 416
12 0 35 0 0 4224 0 73 0 0 0 3
1267 477
1401 477
1401 416
13 0 37 0 0 4224 0 73 0 0 0 3
1267 486
1352 486
1352 418
0 14 39 0 0 4224 0 0 73 0 0 3
1309 417
1309 495
1267 495
7 0 41 0 0 4224 0 74 0 0 0 3
1266 301
1638 301
1638 283
0 8 43 0 0 8320 0 0 74 0 0 3
1591 278
1591 310
1266 310
9 0 45 0 0 4224 0 74 0 0 0 3
1266 319
1548 319
1548 278
10 0 47 0 0 4224 0 74 0 0 0 3
1266 328
1497 328
1497 280
11 0 49 0 0 4224 0 74 0 0 0 3
1266 337
1443 337
1443 280
12 0 51 0 0 4224 0 74 0 0 0 3
1266 346
1397 346
1397 280
13 0 53 0 0 4224 0 74 0 0 0 3
1266 355
1348 355
1348 282
0 14 55 0 0 4224 0 0 74 0 0 3
1303 280
1303 364
1266 364
0 0 3 0 0 4096 0 0 0 127 0 3
1067 476
1067 614
1205 614
0 0 8 0 0 4096 0 0 0 129 0 3
996 200
996 623
1199 623
0 0 4 0 0 8192 0 0 0 128 0 3
949 346
949 485
1198 485
0 0 3 0 0 8192 0 0 0 121 0 4
1032 356
1032 355
1201 355
1201 356
0 0 3 0 0 4096 0 0 0 127 0 3
1032 476
1032 209
1200 209
0 0 2 0 0 8320 0 0 0 123 0 3
937 365
937 218
1200 218
0 0 2 0 0 0 0 0 0 124 0 3
937 494
937 364
1199 364
0 0 2 0 0 0 0 0 0 125 0 4
937 529
937 494
1200 494
1200 493
2 0 2 0 0 0 0 75 0 0 0 4
907 529
937 529
937 632
1199 632
1 0 73 0 0 4224 0 75 0 0 145 3
871 529
74 529
74 474
0 0 3 0 0 8320 0 0 0 213 0 5
84 411
84 397
887 397
887 476
1204 476
0 0 4 0 0 8320 0 0 0 216 0 5
96 367
96 313
949 313
949 346
1205 346
0 0 8 0 0 8320 0 0 0 214 0 5
105 345
105 296
903 296
903 200
1206 200
0 0 5 0 0 4096 0 0 0 131 0 3
1110 448
1110 587
1205 587
0 0 5 0 0 0 0 0 0 132 0 4
1110 318
1110 449
1206 449
1206 448
0 0 5 0 0 8192 0 0 0 133 0 4
1007 173
1110 173
1110 319
1205 319
0 0 5 0 0 8320 0 0 0 218 0 5
225 180
225 60
1007 60
1007 173
1206 173
0 0 6 0 0 4096 0 0 0 135 0 3
1135 440
1135 578
1205 578
0 0 6 0 0 0 0 0 0 136 0 4
1135 309
1135 440
1206 440
1206 439
0 0 6 0 0 8192 0 0 0 137 0 5
1028 164
1135 164
1135 310
1207 310
1207 311
0 0 6 0 0 8320 0 0 0 221 0 5
246 171
246 48
1028 48
1028 164
1206 164
0 0 7 0 0 4096 0 0 0 139 0 3
1160 431
1160 569
1205 569
0 0 7 0 0 0 0 0 0 140 0 4
1159 301
1160 301
1160 431
1204 431
0 0 7 0 0 8192 0 0 0 141 0 5
1049 155
1159 155
1159 301
1207 301
1207 302
0 0 7 0 0 8320 0 0 0 224 0 5
267 162
267 31
1049 31
1049 155
1206 155
0 5 73 0 0 0 0 0 141 145 0 3
173 371
173 216
294 216
0 6 73 0 0 0 0 0 143 144 0 2
173 501
292 501
0 6 73 0 0 0 0 0 142 145 0 3
173 474
173 639
296 639
1 6 73 0 0 0 0 1 144 0 0 4
50 474
173 474
173 371
293 371
0 5 4 0 0 0 0 0 143 216 0 3
137 367
137 492
292 492
0 5 3 0 0 0 0 0 144 213 0 3
153 364
153 362
293 362
0 3 5 0 0 0 0 0 143 217 0 3
225 455
225 456
298 456
1 0 74 0 0 4096 0 76 0 0 236 2
743 567
742 567
1 2 75 0 0 4224 0 77 76 0 0 2
743 533
743 531
1 0 76 0 0 4096 0 78 0 0 237 2
696 566
695 566
1 2 77 0 0 4224 0 79 78 0 0 2
696 532
696 530
1 0 78 0 0 4096 0 80 0 0 228 2
651 567
652 567
1 2 79 0 0 4224 0 81 80 0 0 2
651 533
651 531
1 0 80 0 0 0 0 82 0 0 238 2
601 569
601 569
1 2 81 0 0 4224 0 83 82 0 0 2
601 535
601 533
1 0 82 0 0 0 0 84 0 0 239 2
547 566
547 566
1 2 83 0 0 4224 0 85 84 0 0 2
547 532
547 530
1 0 84 0 0 0 0 86 0 0 240 2
501 567
501 567
1 2 85 0 0 4224 0 87 86 0 0 2
501 533
501 531
1 0 86 0 0 0 0 88 0 0 241 2
452 566
452 566
1 2 87 0 0 4224 0 89 88 0 0 2
452 532
452 530
1 0 88 0 0 0 0 90 0 0 242 2
409 564
409 564
1 2 89 0 0 4224 0 91 90 0 0 2
409 530
409 528
1 0 90 0 0 0 0 92 0 0 243 2
743 430
743 430
1 2 91 0 0 4224 0 93 92 0 0 2
743 396
743 394
1 0 92 0 0 0 0 94 0 0 244 2
696 429
696 429
1 2 93 0 0 4224 0 95 94 0 0 2
696 395
696 393
1 0 94 0 0 0 0 96 0 0 245 2
653 428
653 428
1 2 95 0 0 4224 0 97 96 0 0 2
653 394
653 392
1 0 96 0 0 0 0 98 0 0 246 2
602 430
602 430
1 2 97 0 0 4224 0 99 98 0 0 2
602 396
602 394
1 0 98 0 0 0 0 100 0 0 247 2
548 431
548 431
1 2 99 0 0 4224 0 101 100 0 0 2
548 397
548 395
1 0 100 0 0 0 0 102 0 0 248 2
502 430
502 430
1 2 101 0 0 4224 0 103 102 0 0 2
502 396
502 394
1 0 102 0 0 0 0 104 0 0 249 2
453 430
453 430
1 2 103 0 0 4224 0 105 104 0 0 2
453 396
453 394
1 0 104 0 0 0 0 106 0 0 250 2
410 431
410 431
1 2 105 0 0 4224 0 107 106 0 0 2
410 397
410 395
1 0 106 0 0 0 0 108 0 0 251 2
739 294
739 294
1 2 107 0 0 4224 0 109 108 0 0 2
739 260
739 258
1 0 108 0 0 0 0 110 0 0 252 2
692 292
692 292
1 2 109 0 0 4224 0 111 110 0 0 2
692 258
692 256
1 0 110 0 0 0 0 112 0 0 253 2
649 292
649 292
1 2 111 0 0 4224 0 113 112 0 0 2
649 258
649 256
1 0 112 0 0 0 0 114 0 0 254 2
598 293
598 293
1 2 113 0 0 4224 0 115 114 0 0 2
598 259
598 257
1 0 114 0 0 0 0 116 0 0 255 2
544 291
544 291
1 2 115 0 0 4224 0 117 116 0 0 2
544 257
544 255
1 0 116 0 0 0 0 118 0 0 256 2
498 291
498 291
1 2 117 0 0 4224 0 119 118 0 0 2
498 257
498 255
1 0 118 0 0 0 0 120 0 0 257 2
449 291
449 291
1 2 119 0 0 4224 0 121 120 0 0 2
449 257
449 255
1 0 120 0 0 0 0 122 0 0 258 2
404 289
404 289
1 2 121 0 0 4224 0 123 122 0 0 2
404 255
404 253
1 0 122 0 0 0 0 124 0 0 229 2
740 147
740 147
1 2 123 0 0 4224 0 125 124 0 0 2
740 113
740 111
1 2 124 0 0 4224 0 127 126 0 0 2
693 105
693 103
1 0 125 0 0 0 0 128 0 0 231 2
650 142
650 142
1 2 126 0 0 4224 0 129 128 0 0 2
650 108
650 106
1 0 127 0 0 0 0 130 0 0 232 2
599 144
599 144
1 2 128 0 0 4224 0 131 130 0 0 2
599 110
599 108
1 0 129 0 0 0 0 132 0 0 233 2
545 143
545 143
1 2 130 0 0 4224 0 133 132 0 0 2
545 109
545 107
1 2 131 0 0 4224 0 135 134 0 0 2
499 108
499 106
1 2 132 0 0 4224 0 137 136 0 0 2
450 110
450 108
1 2 133 0 0 4224 0 138 139 0 0 2
404 110
404 108
14 1 134 0 0 8320 0 141 139 0 0 3
370 225
404 225
404 144
0 4 3 0 0 0 0 0 142 212 0 3
153 483
153 621
302 621
0 5 8 0 0 0 0 0 142 214 0 3
123 345
123 630
296 630
0 4 3 0 0 0 0 0 143 213 0 3
153 411
153 483
298 483
1 6 3 0 0 0 0 2 141 0 0 4
52 411
153 411
153 225
294 225
2 4 8 0 0 0 0 140 141 0 0 6
98 346
105 346
105 345
124 345
124 207
300 207
0 1 4 0 0 0 0 0 140 216 0 5
54 367
61 367
61 356
62 356
62 346
1 4 4 0 0 0 0 3 144 0 0 6
55 369
54 369
54 367
138 367
138 353
299 353
0 3 5 0 0 0 0 0 142 218 0 3
225 326
225 594
302 594
0 3 5 0 0 0 0 0 144 225 0 3
225 180
225 326
299 326
0 2 6 0 0 0 0 0 142 220 0 3
246 446
246 585
302 585
0 2 6 0 0 0 0 0 143 221 0 3
246 317
246 447
298 447
0 2 6 0 0 0 0 0 144 226 0 3
246 171
246 317
299 317
0 1 7 0 0 0 0 0 142 223 0 3
267 438
267 576
302 576
0 1 7 0 0 0 0 0 143 224 0 3
267 308
267 438
298 438
0 1 7 0 0 0 0 0 144 227 0 3
267 162
267 308
299 308
1 3 5 0 0 0 0 6 141 0 0 4
75 263
95 263
95 180
300 180
1 2 6 0 0 0 0 5 141 0 0 4
78 214
85 214
85 171
300 171
1 1 7 0 0 0 0 4 141 0 0 3
79 163
79 162
300 162
0 9 78 0 0 8320 0 0 142 0 0 3
652 554
652 594
372 594
7 0 122 0 0 4224 0 141 0 0 0 3
370 162
740 162
740 143
1 8 135 0 0 8320 0 126 141 0 0 3
693 139
693 171
370 171
9 0 125 0 0 4224 0 141 0 0 0 3
370 180
650 180
650 138
10 0 127 0 0 4224 0 141 0 0 0 3
370 189
599 189
599 140
11 0 129 0 0 4224 0 141 0 0 0 3
370 198
545 198
545 140
12 1 136 0 0 4224 0 141 134 0 0 3
370 207
499 207
499 142
13 1 137 0 0 4224 0 141 136 0 0 3
370 216
450 216
450 144
7 0 74 0 0 4224 0 142 0 0 0 3
372 576
742 576
742 557
0 8 76 0 0 8320 0 0 142 0 0 3
695 552
695 585
372 585
10 0 80 0 0 4224 0 142 0 0 0 3
372 603
601 603
601 554
11 0 82 0 0 4224 0 142 0 0 0 3
372 612
547 612
547 554
12 0 84 0 0 4224 0 142 0 0 0 3
372 621
501 621
501 554
13 0 86 0 0 4224 0 142 0 0 0 3
372 630
452 630
452 556
0 14 88 0 0 4224 0 0 142 0 0 3
409 555
409 639
372 639
7 0 90 0 0 4224 0 143 0 0 0 3
368 438
743 438
743 425
0 8 92 0 0 8320 0 0 143 0 0 3
696 420
696 447
368 447
9 0 94 0 0 4224 0 143 0 0 0 3
368 456
653 456
653 420
10 0 96 0 0 4224 0 143 0 0 0 3
368 465
602 465
602 422
11 0 98 0 0 4224 0 143 0 0 0 3
368 474
548 474
548 422
12 0 100 0 0 4224 0 143 0 0 0 3
368 483
502 483
502 422
13 0 102 0 0 4224 0 143 0 0 0 3
368 492
453 492
453 424
0 14 104 0 0 4224 0 0 143 0 0 3
410 423
410 501
368 501
7 0 106 0 0 4224 0 144 0 0 0 3
369 308
739 308
739 289
0 8 108 0 0 8320 0 0 144 0 0 3
692 284
692 317
369 317
9 0 110 0 0 4224 0 144 0 0 0 3
369 326
649 326
649 284
10 0 112 0 0 4224 0 144 0 0 0 3
369 335
598 335
598 286
11 0 114 0 0 4224 0 144 0 0 0 3
369 344
544 344
544 286
12 0 116 0 0 4224 0 144 0 0 0 3
369 353
498 353
498 286
13 0 118 0 0 4224 0 144 0 0 0 3
369 362
449 362
449 288
0 14 120 0 0 4224 0 0 144 0 0 3
404 286
404 371
369 371
7
-27 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
482 769 649 813
497 781 633 811
9 Output 54
-27 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
480 686 693 730
496 697 676 727
12 Input 110110
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
884 536 917 560
892 544 908 560
2 F'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
835 371 864 395
845 379 853 395
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
898 308 927 332
908 316 916 332
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
850 261 887 285
860 269 876 285
2 D'
-27 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 26
479 728 902 772
495 739 885 769
26 F=1, E=1, D=0, IC 7 active
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
