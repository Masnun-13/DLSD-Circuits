CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
52
13 Logic Switch~
5 69 429 0 1 11
0 4
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 S1
-2 -29 12 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3303 0 0
2
5.89953e-315 0
0
13 Logic Switch~
5 98 311 0 1 11
0 5
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 S0
-2 -29 12 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4498 0 0
2
5.89953e-315 0
0
13 Logic Switch~
5 570 720 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9728 0 0
2
5.89953e-315 5.49279e-315
0
13 Logic Switch~
5 564 505 0 1 11
0 36
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3789 0 0
2
5.89953e-315 5.49149e-315
0
13 Logic Switch~
5 575 297 0 1 11
0 42
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3978 0 0
2
5.89953e-315 5.4902e-315
0
13 Logic Switch~
5 566 79 0 1 11
0 48
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3494 0 0
2
5.89953e-315 5.4889e-315
0
13 Logic Switch~
5 571 215 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3507 0 0
2
5.89953e-315 5.48761e-315
0
13 Logic Switch~
5 251 96 0 1 11
0 24
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 B1
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5151 0 0
2
5.89953e-315 5.48631e-315
0
13 Logic Switch~
5 257 323 0 1 11
0 20
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 B2
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3701 0 0
2
5.89953e-315 5.48502e-315
0
13 Logic Switch~
5 285 523 0 1 11
0 16
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 B3
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8585 0 0
2
5.89953e-315 5.48372e-315
0
13 Logic Switch~
5 303 743 0 1 11
0 12
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 B4
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8809 0 0
2
5.89953e-315 5.48243e-315
0
14 Logic Display~
6 907 817 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5993 0 0
2
5.89953e-315 5.48113e-315
0
14 Logic Display~
6 968 728 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8654 0 0
2
5.89953e-315 5.47984e-315
0
9 2-In XOR~
219 802 746 0 3 22
0 28 3 27
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
7223 0 0
2
5.89953e-315 5.47854e-315
0
9 2-In AND~
219 752 844 0 3 22
0 28 3 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3641 0 0
2
5.89953e-315 5.47725e-315
0
8 2-In OR~
219 829 835 0 3 22
0 30 29 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3104 0 0
2
5.89953e-315 5.47595e-315
0
9 2-In AND~
219 648 798 0 3 22
0 31 8 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3296 0 0
2
5.89953e-315 5.47466e-315
0
9 2-In XOR~
219 679 737 0 3 22
0 31 8 28
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8534 0 0
2
5.89953e-315 5.47336e-315
0
14 Logic Display~
6 962 513 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
949 0 0
2
5.89953e-315 5.47207e-315
0
9 2-In XOR~
219 796 531 0 3 22
0 33 2 32
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3371 0 0
2
5.89953e-315 5.47077e-315
0
9 2-In AND~
219 746 630 0 3 22
0 33 2 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7311 0 0
2
5.89953e-315 5.46818e-315
0
8 2-In OR~
219 824 621 0 3 22
0 35 34 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3409 0 0
2
5.89953e-315 5.46559e-315
0
9 2-In AND~
219 642 583 0 3 22
0 36 7 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3526 0 0
2
5.89953e-315 5.463e-315
0
9 2-In XOR~
219 673 522 0 3 22
0 36 7 33
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
4129 0 0
2
5.89953e-315 5.46041e-315
0
14 Logic Display~
6 973 305 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6278 0 0
2
5.89953e-315 5.45782e-315
0
9 2-In XOR~
219 807 323 0 3 22
0 38 6 37
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3482 0 0
2
5.89953e-315 5.45523e-315
0
9 2-In AND~
219 757 421 0 3 22
0 38 6 39
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
8323 0 0
2
5.89953e-315 5.45264e-315
0
8 2-In OR~
219 834 412 0 3 22
0 40 39 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3984 0 0
2
5.89953e-315 5.45005e-315
0
9 2-In AND~
219 653 375 0 3 22
0 42 41 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7622 0 0
2
5.89953e-315 5.44746e-315
0
9 2-In XOR~
219 684 314 0 3 22
0 42 41 38
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
816 0 0
2
5.89953e-315 5.44487e-315
0
9 2-In XOR~
219 675 96 0 3 22
0 48 47 44
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4656 0 0
2
5.89953e-315 5.44228e-315
0
9 2-In AND~
219 644 157 0 3 22
0 48 47 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6356 0 0
2
5.89953e-315 5.43969e-315
0
8 2-In OR~
219 826 197 0 3 22
0 46 45 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7479 0 0
2
5.89953e-315 5.4371e-315
0
9 2-In AND~
219 748 203 0 3 22
0 44 25 45
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
5690 0 0
2
5.89953e-315 5.43451e-315
0
9 2-In XOR~
219 798 105 0 3 22
0 44 25 43
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5617 0 0
2
5.89953e-315 5.43192e-315
0
14 Logic Display~
6 964 87 0 1 2
10 43
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3903 0 0
2
5.89953e-315 5.42933e-315
0
9 Inverter~
13 294 130 0 2 22
0 24 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
4452 0 0
2
5.89953e-315 5.42414e-315
0
9 2-In AND~
219 355 150 0 3 22
0 23 4 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
6282 0 0
2
5.89953e-315 5.41896e-315
0
9 2-In AND~
219 353 53 0 3 22
0 5 24 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
7187 0 0
2
5.89953e-315 5.41378e-315
0
8 2-In OR~
219 426 119 0 3 22
0 21 22 47
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
6866 0 0
2
5.89953e-315 5.4086e-315
0
9 Inverter~
13 300 357 0 2 22
0 20 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
7670 0 0
2
5.89953e-315 5.40342e-315
0
9 2-In AND~
219 361 377 0 3 22
0 19 4 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
951 0 0
2
5.89953e-315 5.39824e-315
0
9 2-In AND~
219 359 280 0 3 22
0 5 20 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
9536 0 0
2
5.89953e-315 5.39306e-315
0
8 2-In OR~
219 433 337 0 3 22
0 17 18 41
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
5495 0 0
2
5.89953e-315 5.38788e-315
0
9 Inverter~
13 328 557 0 2 22
0 16 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
8152 0 0
2
5.89953e-315 5.37752e-315
0
9 2-In AND~
219 389 577 0 3 22
0 15 4 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
6223 0 0
2
5.89953e-315 5.36716e-315
0
9 2-In AND~
219 387 480 0 3 22
0 5 16 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
5441 0 0
2
5.89953e-315 5.3568e-315
0
8 2-In OR~
219 455 545 0 3 22
0 13 14 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U17A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3189 0 0
2
5.89953e-315 5.34643e-315
0
9 Inverter~
13 346 777 0 2 22
0 12 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
8460 0 0
2
5.89953e-315 5.32571e-315
0
9 2-In AND~
219 407 797 0 3 22
0 11 4 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
5179 0 0
2
5.89953e-315 5.30499e-315
0
9 2-In AND~
219 405 700 0 3 22
0 5 12 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
3593 0 0
2
5.89953e-315 5.26354e-315
0
8 2-In OR~
219 471 761 0 3 22
0 9 10 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U17B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
3928 0 0
2
5.89953e-315 0
0
76
0 2 2 0 0 4096 0 0 20 2 0 3
692 638
692 540
780 540
3 2 2 0 0 8320 0 28 21 0 0 7
867 412
867 480
586 480
586 638
692 638
692 639
722 639
0 2 3 0 0 4096 0 0 15 40 0 2
686 853
728 853
0 2 4 0 0 8192 0 0 46 7 0 3
191 588
191 586
365 586
0 2 4 0 0 4096 0 0 38 6 0 3
191 388
191 159
331 159
0 2 4 0 0 0 0 0 42 7 0 3
191 429
191 386
337 386
1 2 4 0 0 8320 0 1 50 0 0 4
81 429
191 429
191 806
383 806
1 0 5 0 0 4096 0 47 0 0 9 2
363 471
145 471
0 1 5 0 0 4224 0 0 51 11 0 3
145 309
145 691
381 691
1 0 5 0 0 0 0 43 0 0 11 2
335 271
145 271
1 1 5 0 0 0 0 39 2 0 0 4
329 44
145 44
145 311
110 311
0 2 6 0 0 4096 0 0 27 59 0 2
692 430
733 430
3 0 7 0 0 4224 0 48 0 0 55 2
488 545
581 545
3 0 8 0 0 8320 0 52 0 0 46 3
504 761
504 760
588 760
3 1 9 0 0 4224 0 51 52 0 0 3
426 700
426 752
458 752
3 2 10 0 0 8320 0 50 52 0 0 3
428 797
428 770
458 770
2 1 11 0 0 8320 0 49 50 0 0 3
367 777
367 788
383 788
1 2 12 0 0 4224 0 11 51 0 0 4
315 743
356 743
356 709
381 709
1 1 12 0 0 0 0 11 49 0 0 3
315 743
315 777
331 777
3 1 13 0 0 4224 0 47 48 0 0 3
408 480
408 536
442 536
3 2 14 0 0 8320 0 46 48 0 0 3
410 577
410 554
442 554
2 1 15 0 0 8320 0 45 46 0 0 3
349 557
349 568
365 568
1 2 16 0 0 4224 0 10 47 0 0 4
297 523
338 523
338 489
363 489
1 1 16 0 0 0 0 10 45 0 0 3
297 523
297 557
313 557
3 1 17 0 0 4224 0 43 44 0 0 3
380 280
380 328
420 328
3 2 18 0 0 8320 0 42 44 0 0 3
382 377
382 346
420 346
2 1 19 0 0 8320 0 41 42 0 0 3
321 357
321 368
337 368
1 2 20 0 0 4224 0 9 43 0 0 4
269 323
310 323
310 289
335 289
1 1 20 0 0 0 0 9 41 0 0 3
269 323
269 357
285 357
3 1 21 0 0 4224 0 39 40 0 0 3
374 53
374 110
413 110
3 2 22 0 0 8320 0 38 40 0 0 3
376 150
376 128
413 128
2 1 23 0 0 8320 0 37 38 0 0 3
315 130
315 141
331 141
1 2 24 0 0 4224 0 8 39 0 0 4
263 96
304 96
304 62
329 62
1 1 24 0 0 0 0 8 37 0 0 3
263 96
263 130
279 130
0 2 25 0 0 4112 0 0 34 69 0 2
682 212
724 212
3 1 26 0 0 4224 0 0 12 37 0 2
884 835
907 835
3 0 26 0 0 0 0 16 0 0 36 2
862 835
885 835
3 1 27 0 0 4224 0 14 13 0 0 2
835 746
968 746
0 1 28 0 0 4096 0 0 14 43 0 2
728 737
786 737
3 2 3 0 0 8320 0 22 14 0 0 7
857 621
857 679
583 679
583 853
687 853
687 755
786 755
3 2 29 0 0 4224 0 15 16 0 0 2
773 844
816 844
3 1 30 0 0 4224 0 17 16 0 0 4
669 798
786 798
786 826
816 826
3 1 28 0 0 8320 0 18 15 0 0 3
712 737
728 737
728 835
0 2 8 0 0 0 0 0 17 46 0 3
604 760
604 807
624 807
0 1 31 0 0 4224 0 0 17 47 0 3
617 720
617 789
624 789
0 2 8 0 0 0 0 0 18 0 0 4
583 760
629 760
629 746
663 746
1 1 31 0 0 0 0 3 18 0 0 4
582 720
629 720
629 728
663 728
3 1 32 0 0 4224 0 20 19 0 0 2
829 531
962 531
0 1 33 0 0 4096 0 0 20 52 0 2
722 522
780 522
3 2 34 0 0 4224 0 21 22 0 0 2
767 630
811 630
3 1 35 0 0 4224 0 23 22 0 0 4
663 583
780 583
780 612
811 612
3 1 33 0 0 8320 0 24 21 0 0 3
706 522
722 522
722 621
0 2 7 0 0 0 0 0 23 55 0 3
598 545
598 592
618 592
0 1 36 0 0 4224 0 0 23 56 0 3
611 505
611 574
618 574
0 2 7 0 0 0 0 0 24 0 0 4
577 545
623 545
623 531
657 531
1 1 36 0 0 0 0 4 24 0 0 4
576 505
623 505
623 513
657 513
3 1 37 0 0 4224 0 26 25 0 0 2
840 323
973 323
0 1 38 0 0 4096 0 0 26 62 0 2
733 314
791 314
3 2 6 0 0 12416 0 33 26 0 0 8
859 197
887 197
887 253
596 253
596 430
692 430
692 332
791 332
3 2 39 0 0 4224 0 27 28 0 0 2
778 421
821 421
3 1 40 0 0 4224 0 29 28 0 0 4
674 375
791 375
791 403
821 403
3 1 38 0 0 8320 0 30 27 0 0 3
717 314
733 314
733 412
0 2 41 0 0 4096 0 0 29 65 0 3
609 337
609 384
629 384
0 1 42 0 0 4224 0 0 29 66 0 3
622 297
622 366
629 366
3 2 41 0 0 4224 0 44 30 0 0 4
466 337
634 337
634 323
668 323
1 1 42 0 0 0 0 5 30 0 0 4
587 297
634 297
634 305
668 305
3 1 43 0 0 4224 0 35 36 0 0 2
831 105
964 105
0 1 44 0 0 4096 0 0 35 72 0 2
724 96
782 96
1 2 25 0 0 8320 0 7 35 0 0 5
583 215
583 212
683 212
683 114
782 114
3 2 45 0 0 12416 0 34 33 0 0 4
769 203
784 203
784 206
813 206
3 1 46 0 0 4224 0 32 33 0 0 4
665 157
782 157
782 188
813 188
3 1 44 0 0 8320 0 31 34 0 0 3
708 96
724 96
724 194
0 2 47 0 0 4096 0 0 32 75 0 3
600 119
600 166
620 166
0 1 48 0 0 4224 0 0 32 76 0 3
613 79
613 148
620 148
3 2 47 0 0 4224 0 40 31 0 0 4
459 119
625 119
625 105
659 105
1 1 48 0 0 0 0 6 31 0 0 4
578 79
625 79
625 87
659 87
65
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
762 840 789 864
767 845 783 861
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
717 856 744 880
722 861 738 877
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
707 818 734 842
712 823 728 839
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
662 776 683 800
668 781 676 797
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
613 808 632 832
618 813 626 829
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
613 761 640 785
618 767 634 783
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
824 745 853 769
830 751 846 767
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
772 758 799 782
777 763 793 779
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
772 708 801 732
778 713 794 729
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
702 715 725 739
709 721 717 737
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
650 695 679 719
656 701 672 717
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
707 289 730 313
714 295 722 311
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
656 273 683 297
661 279 677 295
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
828 322 859 346
835 327 851 343
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
774 284 805 308
781 289 797 305
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
654 748 675 772
660 753 668 769
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
854 813 881 837
859 819 875 835
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
800 849 829 873
806 855 822 871
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
799 802 826 826
804 807 820 823
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
851 598 870 622
856 603 864 619
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
797 634 816 658
802 639 810 655
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
793 587 820 611
798 593 814 609
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
862 390 881 414
867 395 875 411
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
806 427 827 451
812 433 820 449
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
804 380 825 404
810 385 818 401
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
768 420 795 444
773 425 789 441
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
718 434 745 458
723 439 739 455
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
714 393 741 417
719 398 735 414
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
667 353 686 377
672 359 680 375
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
616 385 635 409
621 390 629 406
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
616 338 643 362
621 343 637 359
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
776 335 805 359
782 341 798 357
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
659 325 678 349
664 331 672 347
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
916 828 963 852
923 834 955 850
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
647 481 668 505
653 487 661 503
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
609 546 630 570
615 552 623 568
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
648 533 667 557
653 538 661 554
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
607 593 626 617
612 598 620 614
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
699 498 718 522
704 503 712 519
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
656 561 675 585
661 566 669 582
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
770 492 789 516
775 498 783 514
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
706 599 725 623
711 605 719 621
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
711 641 732 665
717 646 725 662
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
760 625 779 649
765 631 773 647
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
770 543 791 567
776 548 784 564
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
821 530 840 554
826 536 834 552
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
823 104 842 128
828 110 836 126
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
772 117 793 141
778 122 786 138
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
762 199 781 223
767 205 775 221
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
713 215 734 239
719 220 727 236
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
708 173 727 197
713 179 721 195
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
772 66 791 90
777 72 785 88
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
658 135 677 159
663 140 671 156
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
853 172 872 196
858 177 866 193
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
701 72 720 96
706 77 714 93
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
799 208 818 232
804 213 812 229
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
609 167 628 191
614 172 622 188
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
650 107 669 131
655 112 663 128
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
798 161 819 185
804 167 812 183
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
611 120 632 144
617 126 625 142
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
649 55 670 79
655 61 663 77
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
965 111 998 135
973 119 989 135
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
970 330 1003 354
978 338 994 354
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
955 537 988 561
963 545 979 561
2 Y3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
968 752 1001 776
976 760 992 776
2 Y4
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
