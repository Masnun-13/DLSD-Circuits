CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 320 30 200 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 41 513 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 C1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9998 0 0
2
44017.4 0
0
13 Logic Switch~
5 56 385 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-5 -28 9 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3536 0 0
2
44017.4 2
0
13 Logic Switch~
5 59 439 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4597 0 0
2
44017.4 1
0
13 Logic Switch~
5 43 253 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3835 0 0
2
44017.4 0
0
13 Logic Switch~
5 64 145 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
44017.4 0
0
13 Logic Switch~
5 61 91 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-2 -28 5 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
44017.4 0
0
8 2-In OR~
219 265 466 0 3 22
0 8 3 5
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9323 0 0
2
44017.4 0
0
9 2-In AND~
219 179 538 0 3 22
0 6 7 3
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
317 0 0
2
44017.4 7
0
9 Inverter~
13 118 529 0 2 22
0 2 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3108 0 0
2
44017.4 6
0
9 Inverter~
13 86 547 0 2 22
0 4 7
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4299 0 0
2
44017.4 5
0
14 Logic Display~
6 361 448 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
44017.4 3
0
14 Logic Display~
6 366 154 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
44017.4 0
0
8 3-In OR~
219 302 172 0 4 22
0 11 12 10 9
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
6369 0 0
2
44017.4 0
0
9 Inverter~
13 91 253 0 2 22
0 16 15
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9172 0 0
2
44017.4 0
0
9 Inverter~
13 123 235 0 2 22
0 13 14
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7100 0 0
2
44017.4 0
0
9 2-In AND~
219 184 244 0 3 22
0 14 15 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3820 0 0
2
44017.4 0
0
9 2-In AND~
219 222 172 0 3 22
0 17 13 12
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7678 0 0
2
44017.4 0
0
9 2-In AND~
219 161 101 0 3 22
0 18 13 11
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
961 0 0
2
44017.4 0
0
9 Inverter~
13 156 163 0 2 22
0 18 17
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3178 0 0
2
44017.4 0
0
20
1 1 2 0 0 8320 0 3 9 0 0 3
71 439
103 439
103 529
3 2 3 0 0 8320 0 8 7 0 0 4
200 538
235 538
235 475
252 475
1 1 4 0 0 8320 0 1 10 0 0 4
53 513
62 513
62 547
71 547
3 1 5 0 0 4224 0 7 11 0 0 2
298 466
361 466
2 1 6 0 0 4224 0 9 8 0 0 2
139 529
155 529
2 2 7 0 0 4224 0 10 8 0 0 2
107 547
155 547
1 1 8 0 0 16512 0 2 7 0 0 5
68 385
68 386
132 386
132 457
252 457
4 1 9 0 0 4224 0 13 12 0 0 2
335 172
366 172
3 3 10 0 0 4224 0 16 13 0 0 4
205 244
282 244
282 181
289 181
3 1 11 0 0 4224 0 18 13 0 0 4
182 101
264 101
264 163
289 163
3 2 12 0 0 4224 0 17 13 0 0 2
243 172
290 172
1 0 13 0 0 12288 0 15 0 0 18 4
108 235
108 194
81 194
81 145
2 1 14 0 0 4224 0 15 16 0 0 2
144 235
160 235
2 2 15 0 0 4224 0 14 16 0 0 2
112 253
160 253
1 1 16 0 0 4224 0 4 14 0 0 2
55 253
76 253
0 2 13 0 0 8320 0 0 17 18 0 3
97 145
97 181
198 181
1 2 17 0 0 4224 0 17 19 0 0 2
198 163
177 163
1 2 13 0 0 0 0 5 18 0 0 4
76 145
111 145
111 110
137 110
0 1 18 0 0 4224 0 0 19 20 0 3
117 92
117 163
141 163
1 1 18 0 0 0 0 6 18 0 0 3
73 91
73 92
137 92
13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
332 481 407 505
337 485 401 501
8 Y=A+B'C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
22 303 97 347
27 307 91 339
8 Y=A+B'C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
195 510 238 554
200 514 232 546
4 B'C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
133 502 160 526
138 506 154 522
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
88 554 115 578
93 558 109 574
2 C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
332 179 431 203
337 183 425 199
11 AB+A'B+B'C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
93 260 120 284
98 264 114 280
2 C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
138 208 165 232
143 212 159 228
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
200 216 243 260
205 220 237 252
4 B'C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
173 76 200 100
178 80 194 96
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
233 148 268 172
238 152 262 168
3 A'B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
169 132 196 156
174 136 190 152
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
27 9 142 53
32 13 136 45
13 Y=AB+A'B+B'C'
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
