CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
51
13 Logic Switch~
5 562 35 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 S4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3616 0 0
2
5.89957e-315 0
0
13 Logic Switch~
5 483 39 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 S3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5202 0 0
2
5.89957e-315 0
0
13 Logic Switch~
5 518 245 0 1 11
0 17
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 S2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9145 0 0
2
5.89957e-315 0
0
13 Logic Switch~
5 493 252 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 S1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9815 0 0
2
5.89957e-315 0
0
13 Logic Switch~
5 467 253 0 1 11
0 18
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 S0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4766 0 0
2
5.89957e-315 0
0
13 Logic Switch~
5 996 133 0 1 11
0 22
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I31
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8325 0 0
2
5.89957e-315 5.38788e-315
0
13 Logic Switch~
5 974 132 0 1 11
0 21
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I30
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7196 0 0
2
5.89957e-315 5.37752e-315
0
13 Logic Switch~
5 951 131 0 1 11
0 20
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I29
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3567 0 0
2
5.89957e-315 5.36716e-315
0
13 Logic Switch~
5 929 129 0 1 11
0 23
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I28
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5877 0 0
2
5.89957e-315 5.3568e-315
0
13 Logic Switch~
5 910 129 0 1 11
0 24
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I27
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4785 0 0
2
5.89957e-315 5.34643e-315
0
13 Logic Switch~
5 889 129 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I26
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3822 0 0
2
5.89957e-315 5.32571e-315
0
13 Logic Switch~
5 868 129 0 1 11
0 26
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I25
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7640 0 0
2
5.89957e-315 5.30499e-315
0
13 Logic Switch~
5 848 130 0 1 11
0 27
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I24
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9221 0 0
2
5.89957e-315 5.26354e-315
0
13 Logic Switch~
5 809 134 0 1 11
0 30
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I23
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6484 0 0
2
5.89957e-315 5.38788e-315
0
13 Logic Switch~
5 787 133 0 1 11
0 29
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I22
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3689 0 0
2
5.89957e-315 5.37752e-315
0
13 Logic Switch~
5 764 132 0 1 11
0 28
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I21
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3952 0 0
2
5.89957e-315 5.36716e-315
0
13 Logic Switch~
5 742 130 0 1 11
0 31
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I20
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3631 0 0
2
5.89957e-315 5.3568e-315
0
13 Logic Switch~
5 723 130 0 1 11
0 32
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I19
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9359 0 0
2
5.89957e-315 5.34643e-315
0
13 Logic Switch~
5 702 130 0 1 11
0 33
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I18
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5584 0 0
2
5.89957e-315 5.32571e-315
0
13 Logic Switch~
5 681 130 0 1 11
0 34
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I17
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4973 0 0
2
5.89957e-315 5.30499e-315
0
13 Logic Switch~
5 661 131 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I16
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3239 0 0
2
5.89957e-315 5.26354e-315
0
13 Logic Switch~
5 433 132 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I15
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4244 0 0
2
5.89957e-315 5.38788e-315
0
13 Logic Switch~
5 411 131 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I14
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3391 0 0
2
5.89957e-315 5.37752e-315
0
13 Logic Switch~
5 388 130 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I13
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4243 0 0
2
5.89957e-315 5.36716e-315
0
13 Logic Switch~
5 366 128 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3907 0 0
2
5.89957e-315 5.3568e-315
0
13 Logic Switch~
5 347 128 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
728 0 0
2
5.89957e-315 5.34643e-315
0
13 Logic Switch~
5 326 128 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3585 0 0
2
5.89957e-315 5.32571e-315
0
13 Logic Switch~
5 305 128 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3565 0 0
2
5.89957e-315 5.30499e-315
0
13 Logic Switch~
5 285 129 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3966 0 0
2
5.89957e-315 5.26354e-315
0
13 Logic Switch~
5 99 128 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3714 0 0
2
5.89957e-315 5.37752e-315
0
13 Logic Switch~
5 119 127 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3406 0 0
2
5.89957e-315 5.36716e-315
0
13 Logic Switch~
5 140 127 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3132 0 0
2
5.89957e-315 5.3568e-315
0
13 Logic Switch~
5 161 127 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3842 0 0
2
5.89957e-315 5.34643e-315
0
13 Logic Switch~
5 180 127 0 1 11
0 47
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6183 0 0
2
5.89957e-315 5.32571e-315
0
13 Logic Switch~
5 202 129 0 1 11
0 44
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3356 0 0
2
5.89957e-315 5.30499e-315
0
13 Logic Switch~
5 225 130 0 1 11
0 45
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3525 0 0
2
5.89957e-315 5.26354e-315
0
13 Logic Switch~
5 247 131 0 1 11
0 46
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3800 0 0
2
5.89957e-315 0
0
14 Logic Display~
6 594 446 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
346 0 0
2
5.89957e-315 0
0
9 Inverter~
13 585 76 0 2 22
0 9 7
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U8B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
3169 0 0
2
5.89957e-315 0
0
9 Inverter~
13 502 74 0 2 22
0 10 8
0
0 0 608 270
5 74F04
-18 -19 17 -11
3 U8A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
4826 0 0
2
5.89957e-315 0
0
8 2-In OR~
219 585 131 0 3 22
0 7 8 3
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U7A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3971 0 0
2
5.89957e-315 0
0
8 2-In OR~
219 546 131 0 3 22
0 7 10 4
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U5D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3607 0 0
2
5.89957e-315 0
0
8 2-In OR~
219 506 131 0 3 22
0 9 8 5
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U5C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3506 0 0
2
5.89957e-315 0
0
8 2-In OR~
219 468 130 0 3 22
0 9 10 6
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U5B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7829 0 0
2
5.89957e-315 0
0
8 2-In OR~
219 496 442 0 3 22
0 11 12 2
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U5A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3890 0 0
2
5.89957e-315 0
0
8 2-In OR~
219 819 347 0 3 22
0 14 15 11
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U6B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3126 0 0
2
5.89957e-315 0
0
8 2-In OR~
219 229 344 0 3 22
0 16 13 12
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U6A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3935 0 0
2
5.89957e-315 0
0
7 74LS151
20 901 238 0 14 29
0 22 21 20 23 24 25 26 27 3
17 19 18 14 52
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U4
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
9746 0 0
2
5.89957e-315 0
0
7 74LS151
20 714 235 0 14 29
0 30 29 28 31 32 33 34 35 4
17 19 18 15 53
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U3
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7330 0 0
2
5.89957e-315 0
0
7 74LS151
20 338 237 0 14 29
0 38 37 36 39 40 41 42 43 5
17 19 18 16 54
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U2
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3972 0 0
2
5.89957e-315 0
0
7 74LS151
20 152 237 0 14 29
0 46 45 44 47 48 49 50 51 6
17 19 18 13 55
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U1
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7818 0 0
2
5.89957e-315 5.38788e-315
0
65
3 1 2 0 0 8320 0 45 38 0 0 4
499 472
499 486
594 486
594 464
3 9 3 0 0 8320 0 41 48 0 0 4
588 161
588 375
927 375
927 271
3 9 4 0 0 8320 0 42 49 0 0 4
549 161
549 333
740 333
740 268
3 9 5 0 0 4224 0 43 50 0 0 4
509 161
509 328
364 328
364 270
3 9 6 0 0 8320 0 44 51 0 0 4
471 160
471 312
178 312
178 270
2 1 7 0 0 8192 0 39 41 0 0 3
588 94
597 94
597 115
2 1 7 0 0 4224 0 39 42 0 0 3
588 94
558 94
558 115
0 2 8 0 0 4224 0 0 41 9 0 3
505 108
579 108
579 115
2 2 8 0 0 0 0 40 43 0 0 4
505 92
505 108
500 108
500 115
1 0 9 0 0 4096 0 39 0 0 13 2
588 58
562 58
1 0 10 0 0 4096 0 40 0 0 14 2
505 56
505 51
1 0 9 0 0 4096 0 43 0 0 13 2
518 115
518 78
1 1 9 0 0 8320 0 1 44 0 0 4
562 47
562 78
480 78
480 114
1 2 10 0 0 8320 0 2 42 0 0 3
483 51
540 51
540 115
2 1 10 0 0 0 0 44 2 0 0 3
462 114
462 51
483 51
3 1 11 0 0 8320 0 46 45 0 0 4
822 377
822 416
508 416
508 426
3 2 12 0 0 8320 0 47 45 0 0 4
232 374
232 415
490 415
490 426
13 2 13 0 0 8320 0 51 47 0 0 4
124 264
124 322
223 322
223 328
1 13 14 0 0 12416 0 46 48 0 0 4
831 331
831 318
873 318
873 265
2 13 15 0 0 8320 0 46 49 0 0 4
813 331
813 316
686 316
686 262
1 13 16 0 0 8320 0 47 50 0 0 4
241 328
241 318
310 318
310 264
10 0 17 0 0 4096 0 50 0 0 25 2
355 264
355 298
10 0 17 0 0 4096 0 49 0 0 24 2
731 262
731 298
0 10 17 0 0 4224 0 0 48 25 0 3
518 298
918 298
918 265
1 10 17 0 0 0 0 3 51 0 0 4
518 257
518 298
169 298
169 264
12 0 18 0 0 4096 0 49 0 0 31 2
713 262
713 276
11 0 19 0 0 4096 0 49 0 0 28 2
722 262
722 287
0 11 19 0 0 4224 0 0 48 30 0 3
493 287
909 287
909 265
11 0 19 0 0 0 0 50 0 0 30 2
346 264
346 287
1 11 19 0 0 0 0 4 51 0 0 4
493 264
493 287
160 287
160 264
0 12 18 0 0 4224 0 0 48 33 0 3
467 276
900 276
900 265
0 12 18 0 0 0 0 0 51 33 0 3
337 276
151 276
151 264
12 1 18 0 0 0 0 50 5 0 0 4
337 264
337 276
467 276
467 265
1 3 20 0 0 8320 0 8 48 0 0 4
951 143
951 182
909 182
909 201
1 2 21 0 0 8320 0 7 48 0 0 4
974 144
974 191
918 191
918 201
1 1 22 0 0 8320 0 48 6 0 0 4
927 201
927 197
996 197
996 145
4 1 23 0 0 20608 0 48 9 0 0 6
900 201
900 194
905 194
905 178
929 178
929 141
1 5 24 0 0 4224 0 10 48 0 0 6
910 141
910 171
902 171
902 187
891 187
891 201
1 6 25 0 0 4224 0 11 48 0 0 4
889 141
889 180
882 180
882 201
7 1 26 0 0 4224 0 48 12 0 0 3
873 201
873 141
868 141
1 8 27 0 0 4224 0 13 48 0 0 4
848 142
848 194
864 194
864 201
1 3 28 0 0 8320 0 16 49 0 0 4
764 144
764 183
722 183
722 198
1 2 29 0 0 8320 0 15 49 0 0 4
787 145
787 192
731 192
731 198
1 1 30 0 0 4224 0 49 14 0 0 3
740 198
809 198
809 146
4 1 31 0 0 20608 0 49 17 0 0 6
713 198
713 195
718 195
718 179
742 179
742 142
1 5 32 0 0 4224 0 18 49 0 0 6
723 142
723 172
715 172
715 188
704 188
704 198
1 6 33 0 0 4224 0 19 49 0 0 4
702 142
702 181
695 181
695 198
7 1 34 0 0 4224 0 49 20 0 0 3
686 198
686 142
681 142
1 8 35 0 0 4224 0 21 49 0 0 4
661 143
661 195
677 195
677 198
1 3 36 0 0 8320 0 24 50 0 0 4
388 142
388 181
346 181
346 200
1 2 37 0 0 8320 0 23 50 0 0 4
411 143
411 190
355 190
355 200
1 1 38 0 0 8320 0 50 22 0 0 4
364 200
364 196
433 196
433 144
4 1 39 0 0 20608 0 50 25 0 0 6
337 200
337 193
342 193
342 177
366 177
366 140
1 5 40 0 0 4224 0 26 50 0 0 6
347 140
347 170
339 170
339 186
328 186
328 200
1 6 41 0 0 4224 0 27 50 0 0 4
326 140
326 179
319 179
319 200
7 1 42 0 0 4224 0 50 28 0 0 3
310 200
310 140
305 140
1 8 43 0 0 4224 0 29 50 0 0 4
285 141
285 193
301 193
301 200
1 3 44 0 0 8320 0 35 51 0 0 4
202 141
202 180
160 180
160 200
1 2 45 0 0 8320 0 36 51 0 0 4
225 142
225 189
169 189
169 200
1 1 46 0 0 8320 0 51 37 0 0 4
178 200
178 195
247 195
247 143
4 1 47 0 0 20608 0 51 34 0 0 6
151 200
151 192
156 192
156 176
180 176
180 139
1 5 48 0 0 4224 0 33 51 0 0 6
161 139
161 169
153 169
153 185
142 185
142 200
1 6 49 0 0 4224 0 32 51 0 0 4
140 139
140 178
133 178
133 200
7 1 50 0 0 4224 0 51 31 0 0 3
124 200
124 139
119 139
1 8 51 0 0 4224 0 30 51 0 0 4
99 140
99 192
115 192
115 200
1
-19 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 63
74 422 335 505
83 428 325 491
63 Input: 11010 = 26
S3=1 S4=1 IC4 active
Output I26=1, verified
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
