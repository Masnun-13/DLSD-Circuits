CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
89
13 Logic Switch~
5 1269 251 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 S7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4389 0 0
2
44111.4 0
0
13 Logic Switch~
5 1210 230 0 1 11
0 3
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 S6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7762 0 0
2
44111.4 1
0
13 Logic Switch~
5 1270 395 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 S5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6723 0 0
2
44111.4 2
0
13 Logic Switch~
5 1227 386 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 S4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6871 0 0
2
44111.4 3
0
13 Logic Switch~
5 1184 376 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 S3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4198 0 0
2
44111.4 4
0
13 Logic Switch~
5 585 174 0 10 11
0 58 0 0 0 0 0 0 0 0
1
0
0 0 21344 180
2 5V
-7 -16 7 -8
2 S2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
970 0 0
2
44111.4 5
0
13 Logic Switch~
5 551 105 0 1 11
0 59
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 S0
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
319 0 0
2
44111.4 6
0
13 Logic Switch~
5 576 135 0 1 11
0 60
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 S1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3663 0 0
2
44111.4 7
0
13 Logic Switch~
5 89 446 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I32
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3512 0 0
2
5.89957e-315 0
0
13 Logic Switch~
5 109 445 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I33
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7555 0 0
2
5.89957e-315 5.26354e-315
0
13 Logic Switch~
5 130 445 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I34
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9776 0 0
2
5.89957e-315 5.30499e-315
0
13 Logic Switch~
5 151 445 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I35
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6596 0 0
2
5.89957e-315 5.32571e-315
0
13 Logic Switch~
5 170 445 0 1 11
0 21
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I36
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6750 0 0
2
5.89957e-315 5.34643e-315
0
13 Logic Switch~
5 192 447 0 1 11
0 18
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I37
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9636 0 0
2
5.89957e-315 5.3568e-315
0
13 Logic Switch~
5 215 448 0 1 11
0 19
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I38
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5369 0 0
2
5.89957e-315 5.36716e-315
0
13 Logic Switch~
5 237 449 0 1 11
0 20
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I39
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8555 0 0
2
5.89957e-315 5.37752e-315
0
13 Logic Switch~
5 986 447 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I63
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4690 0 0
2
5.89957e-315 5.38788e-315
0
13 Logic Switch~
5 964 446 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I62
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9145 0 0
2
5.89957e-315 5.39306e-315
0
13 Logic Switch~
5 941 445 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I61
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5246 0 0
2
5.89957e-315 5.39824e-315
0
13 Logic Switch~
5 919 443 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I60
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9111 0 0
2
5.89957e-315 5.40342e-315
0
13 Logic Switch~
5 900 443 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I59
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6717 0 0
2
5.89957e-315 5.4086e-315
0
13 Logic Switch~
5 879 443 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I58
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3487 0 0
2
5.89957e-315 5.41378e-315
0
13 Logic Switch~
5 858 443 0 1 11
0 32
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I57
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9604 0 0
2
5.89957e-315 5.41896e-315
0
13 Logic Switch~
5 838 444 0 1 11
0 33
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I56
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3921 0 0
2
5.89957e-315 5.42414e-315
0
13 Logic Switch~
5 799 447 0 1 11
0 36
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I55
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8146 0 0
2
5.89957e-315 5.42933e-315
0
13 Logic Switch~
5 777 446 0 1 11
0 35
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I54
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4506 0 0
2
5.89957e-315 5.43192e-315
0
13 Logic Switch~
5 754 445 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I53
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5386 0 0
2
5.89957e-315 5.43451e-315
0
13 Logic Switch~
5 732 443 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I52
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7847 0 0
2
5.89957e-315 5.4371e-315
0
13 Logic Switch~
5 713 443 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I51
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9261 0 0
2
5.89957e-315 5.43969e-315
0
13 Logic Switch~
5 692 443 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I50
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8231 0 0
2
5.89957e-315 5.44228e-315
0
13 Logic Switch~
5 671 443 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I49
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3756 0 0
2
5.89957e-315 5.44487e-315
0
13 Logic Switch~
5 651 444 0 1 11
0 41
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I48
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6760 0 0
2
5.89957e-315 5.44746e-315
0
13 Logic Switch~
5 423 449 0 1 11
0 44
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I47
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
351 0 0
2
5.89957e-315 5.45005e-315
0
13 Logic Switch~
5 401 448 0 1 11
0 43
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I46
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5352 0 0
2
5.89957e-315 5.45264e-315
0
13 Logic Switch~
5 378 447 0 1 11
0 42
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I45
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
485 0 0
2
5.89957e-315 5.45523e-315
0
13 Logic Switch~
5 356 445 0 1 11
0 45
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I44
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
452 0 0
2
5.89957e-315 5.45782e-315
0
13 Logic Switch~
5 337 445 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I43
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
643 0 0
2
5.89957e-315 5.46041e-315
0
13 Logic Switch~
5 316 445 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I42
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5563 0 0
2
5.89957e-315 5.463e-315
0
13 Logic Switch~
5 295 445 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I41
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
934 0 0
2
5.89957e-315 5.46559e-315
0
13 Logic Switch~
5 275 446 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I40
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3240 0 0
2
5.89957e-315 5.46818e-315
0
13 Logic Switch~
5 996 133 0 1 11
0 67
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I31
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3233 0 0
2
5.89957e-315 5.47077e-315
0
13 Logic Switch~
5 974 132 0 1 11
0 66
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I30
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3635 0 0
2
5.89957e-315 5.47207e-315
0
13 Logic Switch~
5 951 131 0 1 11
0 65
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I29
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3547 0 0
2
5.89957e-315 5.47336e-315
0
13 Logic Switch~
5 929 129 0 1 11
0 68
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I28
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
483 0 0
2
5.89957e-315 5.47466e-315
0
13 Logic Switch~
5 910 129 0 1 11
0 69
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I27
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6126 0 0
2
5.89957e-315 5.47595e-315
0
13 Logic Switch~
5 889 129 0 1 11
0 70
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I26
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7368 0 0
2
5.89957e-315 5.47725e-315
0
13 Logic Switch~
5 868 129 0 1 11
0 71
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I25
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3925 0 0
2
5.89957e-315 5.47854e-315
0
13 Logic Switch~
5 848 130 0 1 11
0 72
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I24
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6187 0 0
2
5.89957e-315 5.47984e-315
0
13 Logic Switch~
5 809 134 0 1 11
0 75
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I23
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5866 0 0
2
5.89957e-315 5.48113e-315
0
13 Logic Switch~
5 787 133 0 1 11
0 74
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I22
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6650 0 0
2
5.89957e-315 5.48243e-315
0
13 Logic Switch~
5 764 132 0 1 11
0 73
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I21
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8814 0 0
2
5.89957e-315 5.48372e-315
0
13 Logic Switch~
5 742 130 0 1 11
0 76
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I20
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4714 0 0
2
5.89957e-315 5.48502e-315
0
13 Logic Switch~
5 723 130 0 1 11
0 77
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I19
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9875 0 0
2
5.89957e-315 5.48631e-315
0
13 Logic Switch~
5 702 130 0 1 11
0 78
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I18
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8220 0 0
2
5.89957e-315 5.48761e-315
0
13 Logic Switch~
5 681 130 0 1 11
0 79
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 I17
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3691 0 0
2
5.89957e-315 5.4889e-315
0
13 Logic Switch~
5 661 131 0 10 11
0 80 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I16
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5196 0 0
2
5.89957e-315 5.4902e-315
0
13 Logic Switch~
5 433 132 0 10 11
0 83 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I15
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6182 0 0
2
5.89957e-315 5.49149e-315
0
13 Logic Switch~
5 411 131 0 10 11
0 82 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I14
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6326 0 0
2
5.89957e-315 5.49279e-315
0
13 Logic Switch~
5 388 130 0 10 11
0 81 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I13
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3247 0 0
2
5.89957e-315 5.49408e-315
0
13 Logic Switch~
5 366 128 0 10 11
0 84 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5235 0 0
2
5.89957e-315 5.49538e-315
0
13 Logic Switch~
5 347 128 0 10 11
0 85 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9260 0 0
2
5.89957e-315 5.49667e-315
0
13 Logic Switch~
5 326 128 0 10 11
0 86 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 I10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
583 0 0
2
5.89957e-315 5.49797e-315
0
13 Logic Switch~
5 305 128 0 10 11
0 87 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3471 0 0
2
5.89957e-315 5.49926e-315
0
13 Logic Switch~
5 285 129 0 10 11
0 88 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7124 0 0
2
5.89957e-315 5.50056e-315
0
13 Logic Switch~
5 99 128 0 10 11
0 96 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6160 0 0
2
5.89957e-315 5.50185e-315
0
13 Logic Switch~
5 119 127 0 10 11
0 95 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4732 0 0
2
5.89957e-315 5.50315e-315
0
13 Logic Switch~
5 140 127 0 10 11
0 94 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8836 0 0
2
5.89957e-315 5.50444e-315
0
13 Logic Switch~
5 161 127 0 10 11
0 93 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3346 0 0
2
5.89957e-315 5.50574e-315
0
13 Logic Switch~
5 180 127 0 10 11
0 92 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8546 0 0
2
5.89957e-315 5.50703e-315
0
13 Logic Switch~
5 202 129 0 10 11
0 89 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8607 0 0
2
5.89957e-315 5.50833e-315
0
13 Logic Switch~
5 225 130 0 10 11
0 90 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 I6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5781 0 0
2
5.89957e-315 5.50963e-315
0
13 Logic Switch~
5 247 131 0 1 11
0 91
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 I7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6991 0 0
2
5.89957e-315 5.51092e-315
0
14 Logic Display~
6 722 746 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9631 0 0
2
44111.4 8
0
7 74LS138
19 1109 376 0 14 29
0 13 14 15 4 3 3 6 5 7
8 9 10 11 12
0
0 0 5088 180
7 74LS138
-25 -62 24 -54
3 U13
-11 -72 10 -64
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8381 0 0
2
44111.4 9
0
7 74LS151
20 142 548 0 14 29
0 20 19 18 21 22 23 24 25 8
58 60 59 54 97
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U7
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
6697 0 0
2
5.89957e-315 5.51222e-315
0
7 74LS151
20 891 552 0 14 29
0 28 27 26 29 30 31 32 33 6
58 60 59 55 98
0
0 0 4832 270
6 74F151
-21 -60 21 -52
3 U11
52 -10 73 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3463 0 0
2
5.89957e-315 5.51286e-315
0
7 74LS151
20 704 550 0 14 29
0 36 35 34 37 38 39 40 41 5
58 60 59 56 99
0
0 0 4832 270
6 74F151
-21 -60 21 -52
3 U10
52 -10 73 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
9605 0 0
2
5.89957e-315 5.51351e-315
0
7 74LS151
20 328 548 0 14 29
0 44 43 42 45 46 47 48 49 7
58 60 59 57 100
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U8
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
936 0 0
2
5.89957e-315 5.51416e-315
0
8 2-In OR~
219 494 771 0 3 22
0 50 51 2
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U5A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9813 0 0
2
5.89957e-315 5.51481e-315
0
8 2-In OR~
219 612 723 0 3 22
0 53 101 50
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U9D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 6 0
1 U
5286 0 0
2
5.89957e-315 5.51545e-315
0
8 2-In OR~
219 398 669 0 3 22
0 16 17 51
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U9C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
9179 0 0
2
5.89957e-315 5.5161e-315
0
8 2-In OR~
219 219 658 0 3 22
0 57 54 52
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U9B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3718 0 0
2
5.89957e-315 5.51675e-315
0
8 2-In OR~
219 809 661 0 3 22
0 55 56 53
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U9A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4375 0 0
2
5.89957e-315 5.5174e-315
0
8 2-In OR~
219 819 347 0 3 22
0 62 63 16
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U6B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3616 0 0
2
5.89957e-315 5.51804e-315
0
8 2-In OR~
219 229 344 0 3 22
0 64 61 17
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U6A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7808 0 0
2
5.89957e-315 5.51869e-315
0
7 74LS151
20 901 238 0 14 29
0 67 66 65 68 69 70 71 72 9
58 60 59 62 102
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U4
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7498 0 0
2
5.89957e-315 5.51934e-315
0
7 74LS151
20 714 235 0 14 29
0 75 74 73 76 77 78 79 80 10
58 60 59 63 103
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U3
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
9736 0 0
2
5.89957e-315 5.51999e-315
0
7 74LS151
20 338 237 0 14 29
0 83 82 81 84 85 86 87 88 11
58 60 59 64 104
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U2
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
9454 0 0
2
5.89957e-315 5.52063e-315
0
7 74LS151
20 152 237 0 14 29
0 91 90 89 92 93 94 95 96 12
58 60 59 61 105
0
0 0 4832 270
6 74F151
-21 -60 21 -52
2 U1
55 -10 69 -2
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
4639 0 0
2
5.89957e-315 5.52128e-315
0
117
3 1 2 0 0 4224 0 79 73 0 0 3
497 801
722 801
722 764
5 0 3 0 0 8192 0 74 0 0 3 3
1147 341
1155 341
1155 332
1 6 3 0 0 8320 0 2 74 0 0 4
1196 230
1172 230
1172 332
1147 332
4 1 4 0 0 16512 0 74 1 0 0 6
1141 350
1162 350
1162 341
1245 341
1245 251
1255 251
8 9 5 0 0 12416 0 74 77 0 0 5
1071 386
1049 386
1049 619
730 619
730 583
9 7 6 0 0 8320 0 76 74 0 0 4
917 585
1061 585
1061 395
1071 395
9 9 7 0 0 8320 0 78 74 0 0 5
354 581
354 641
1040 641
1040 377
1071 377
10 9 8 0 0 12416 0 74 75 0 0 5
1071 368
1025 368
1025 625
168 625
168 581
9 11 9 0 0 8320 0 86 74 0 0 3
927 271
927 359
1071 359
12 9 10 0 0 4224 0 74 87 0 0 3
1071 350
740 350
740 268
9 13 11 0 0 8320 0 88 74 0 0 3
364 270
364 341
1071 341
9 14 12 0 0 8320 0 89 74 0 0 3
178 270
178 332
1071 332
1 1 13 0 0 4224 0 74 3 0 0 2
1141 395
1256 395
2 1 14 0 0 4224 0 74 4 0 0 2
1141 386
1213 386
3 1 15 0 0 8320 0 74 5 0 0 3
1141 377
1141 376
1170 376
3 1 16 0 0 4224 0 84 81 0 0 3
822 377
410 377
410 653
2 3 17 0 0 4224 0 81 85 0 0 4
392 653
392 386
232 386
232 374
1 3 18 0 0 8320 0 14 75 0 0 4
192 459
192 498
150 498
150 511
1 2 19 0 0 8320 0 15 75 0 0 4
215 460
215 507
159 507
159 511
1 1 20 0 0 8320 0 75 16 0 0 4
168 511
168 513
237 513
237 461
4 1 21 0 0 20608 0 75 13 0 0 6
141 511
141 510
146 510
146 494
170 494
170 457
1 5 22 0 0 4224 0 12 75 0 0 6
151 457
151 487
143 487
143 503
132 503
132 511
1 6 23 0 0 4224 0 11 75 0 0 4
130 457
130 496
123 496
123 511
7 1 24 0 0 4224 0 75 10 0 0 3
114 511
114 457
109 457
1 8 25 0 0 4224 0 9 75 0 0 4
89 458
89 510
105 510
105 511
1 3 26 0 0 8320 0 19 76 0 0 4
941 457
941 496
899 496
899 515
1 2 27 0 0 8320 0 18 76 0 0 4
964 458
964 505
908 505
908 515
1 1 28 0 0 8320 0 76 17 0 0 4
917 515
917 511
986 511
986 459
4 1 29 0 0 20608 0 76 20 0 0 6
890 515
890 508
895 508
895 492
919 492
919 455
1 5 30 0 0 4224 0 21 76 0 0 6
900 455
900 485
892 485
892 501
881 501
881 515
1 6 31 0 0 4224 0 22 76 0 0 4
879 455
879 494
872 494
872 515
7 1 32 0 0 4224 0 76 23 0 0 3
863 515
863 455
858 455
1 8 33 0 0 4224 0 24 76 0 0 4
838 456
838 508
854 508
854 515
1 3 34 0 0 8320 0 27 77 0 0 4
754 457
754 496
712 496
712 513
1 2 35 0 0 8320 0 26 77 0 0 4
777 458
777 505
721 505
721 513
1 1 36 0 0 8320 0 77 25 0 0 4
730 513
730 511
799 511
799 459
4 1 37 0 0 20608 0 77 28 0 0 6
703 513
703 508
708 508
708 492
732 492
732 455
1 5 38 0 0 4224 0 29 77 0 0 6
713 455
713 485
705 485
705 501
694 501
694 513
1 6 39 0 0 4224 0 30 77 0 0 4
692 455
692 494
685 494
685 513
7 1 40 0 0 4224 0 77 31 0 0 3
676 513
676 455
671 455
1 8 41 0 0 4224 0 32 77 0 0 4
651 456
651 508
667 508
667 513
1 3 42 0 0 8320 0 35 78 0 0 4
378 459
378 498
336 498
336 511
1 2 43 0 0 8320 0 34 78 0 0 4
401 460
401 507
345 507
345 511
1 1 44 0 0 8320 0 78 33 0 0 4
354 511
354 513
423 513
423 461
4 1 45 0 0 20608 0 78 36 0 0 6
327 511
327 510
332 510
332 494
356 494
356 457
1 5 46 0 0 4224 0 37 78 0 0 6
337 457
337 487
329 487
329 503
318 503
318 511
1 6 47 0 0 4224 0 38 78 0 0 4
316 457
316 496
309 496
309 511
7 1 48 0 0 4224 0 78 39 0 0 3
300 511
300 457
295 457
1 8 49 0 0 4224 0 40 78 0 0 4
275 458
275 510
291 510
291 511
3 1 50 0 0 4224 0 80 79 0 0 3
615 753
506 753
506 755
3 2 51 0 0 8320 0 81 79 0 0 4
401 699
401 753
488 753
488 755
0 3 52 0 0 8320 0 0 82 0 0 4
604 713
604 699
222 699
222 688
3 1 53 0 0 8320 0 83 80 0 0 4
812 691
812 699
624 699
624 707
13 2 54 0 0 8320 0 75 82 0 0 4
114 575
114 636
213 636
213 642
1 13 55 0 0 12416 0 83 76 0 0 4
821 645
821 632
863 632
863 579
2 13 56 0 0 8320 0 83 77 0 0 4
803 645
803 630
676 630
676 577
1 13 57 0 0 8320 0 82 78 0 0 4
231 642
231 632
300 632
300 575
10 0 58 0 0 4096 0 78 0 0 61 2
345 575
345 612
10 0 58 0 0 0 0 77 0 0 60 2
721 577
721 612
0 10 58 0 0 4224 0 0 76 61 0 3
508 612
908 612
908 579
0 10 58 0 0 0 0 0 75 77 0 4
508 298
508 612
159 612
159 575
12 0 59 0 0 4096 0 77 0 0 67 2
703 577
703 593
11 0 60 0 0 4096 0 77 0 0 64 2
712 577
712 601
0 11 60 0 0 4224 0 0 76 66 0 3
483 601
899 601
899 579
11 0 60 0 0 0 0 78 0 0 66 2
336 575
336 601
0 11 60 0 0 0 0 0 75 82 0 4
483 287
483 601
150 601
150 575
0 12 59 0 0 8320 0 0 76 69 0 4
457 590
457 593
890 593
890 579
0 12 59 0 0 0 0 0 75 69 0 3
327 590
141 590
141 575
12 0 59 0 0 0 0 78 0 0 85 4
327 575
327 590
457 590
457 276
13 2 61 0 0 8320 0 89 85 0 0 4
124 264
124 322
223 322
223 328
1 13 62 0 0 12416 0 84 86 0 0 4
831 331
831 318
873 318
873 265
2 13 63 0 0 8320 0 84 87 0 0 4
813 331
813 316
686 316
686 262
1 13 64 0 0 8320 0 85 88 0 0 4
241 328
241 318
310 318
310 264
10 0 58 0 0 0 0 88 0 0 77 2
355 264
355 298
10 0 58 0 0 0 0 87 0 0 76 2
731 262
731 298
0 10 58 0 0 0 0 0 86 77 0 3
518 298
918 298
918 265
1 10 58 0 0 0 0 6 89 0 0 5
571 174
518 174
518 298
169 298
169 264
12 0 59 0 0 0 0 87 0 0 83 2
713 262
713 276
11 0 60 0 0 0 0 87 0 0 80 2
722 262
722 287
0 11 60 0 0 0 0 0 86 82 0 3
493 287
909 287
909 265
11 0 60 0 0 0 0 88 0 0 82 2
346 264
346 287
1 11 60 0 0 0 0 8 89 0 0 5
562 135
493 135
493 287
160 287
160 264
0 12 59 0 0 0 0 0 86 85 0 3
467 276
900 276
900 265
0 12 59 0 0 0 0 0 89 85 0 3
337 276
151 276
151 264
12 1 59 0 0 0 0 88 7 0 0 5
337 264
337 276
467 276
467 105
537 105
1 3 65 0 0 8320 0 43 86 0 0 4
951 143
951 182
909 182
909 201
1 2 66 0 0 8320 0 42 86 0 0 4
974 144
974 191
918 191
918 201
1 1 67 0 0 8320 0 86 41 0 0 4
927 201
927 197
996 197
996 145
4 1 68 0 0 20608 0 86 44 0 0 6
900 201
900 194
905 194
905 178
929 178
929 141
1 5 69 0 0 4224 0 45 86 0 0 6
910 141
910 171
902 171
902 187
891 187
891 201
1 6 70 0 0 4224 0 46 86 0 0 4
889 141
889 180
882 180
882 201
7 1 71 0 0 4224 0 86 47 0 0 3
873 201
873 141
868 141
1 8 72 0 0 4224 0 48 86 0 0 4
848 142
848 194
864 194
864 201
1 3 73 0 0 8320 0 51 87 0 0 4
764 144
764 183
722 183
722 198
1 2 74 0 0 8320 0 50 87 0 0 4
787 145
787 192
731 192
731 198
1 1 75 0 0 4224 0 87 49 0 0 3
740 198
809 198
809 146
4 1 76 0 0 20608 0 87 52 0 0 6
713 198
713 195
718 195
718 179
742 179
742 142
1 5 77 0 0 4224 0 53 87 0 0 6
723 142
723 172
715 172
715 188
704 188
704 198
1 6 78 0 0 4224 0 54 87 0 0 4
702 142
702 181
695 181
695 198
7 1 79 0 0 4224 0 87 55 0 0 3
686 198
686 142
681 142
1 8 80 0 0 4224 0 56 87 0 0 4
661 143
661 195
677 195
677 198
1 3 81 0 0 8320 0 59 88 0 0 4
388 142
388 181
346 181
346 200
1 2 82 0 0 8320 0 58 88 0 0 4
411 143
411 190
355 190
355 200
1 1 83 0 0 8320 0 88 57 0 0 4
364 200
364 196
433 196
433 144
4 1 84 0 0 20608 0 88 60 0 0 6
337 200
337 193
342 193
342 177
366 177
366 140
1 5 85 0 0 4224 0 61 88 0 0 6
347 140
347 170
339 170
339 186
328 186
328 200
1 6 86 0 0 4224 0 62 88 0 0 4
326 140
326 179
319 179
319 200
7 1 87 0 0 4224 0 88 63 0 0 3
310 200
310 140
305 140
1 8 88 0 0 4224 0 64 88 0 0 4
285 141
285 193
301 193
301 200
1 3 89 0 0 8320 0 70 89 0 0 4
202 141
202 180
160 180
160 200
1 2 90 0 0 8320 0 71 89 0 0 4
225 142
225 189
169 189
169 200
1 1 91 0 0 8320 0 89 72 0 0 4
178 200
178 195
247 195
247 143
4 1 92 0 0 20608 0 89 69 0 0 6
151 200
151 192
156 192
156 176
180 176
180 139
1 5 93 0 0 4224 0 68 89 0 0 6
161 139
161 169
153 169
153 185
142 185
142 200
1 6 94 0 0 4224 0 67 89 0 0 4
140 139
140 178
133 178
133 200
7 1 95 0 0 4224 0 89 66 0 0 3
124 200
124 139
119 139
1 8 96 0 0 4224 0 65 89 0 0 4
99 140
99 192
115 192
115 200
1
-19 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 69
960 656 1271 739
972 666 1258 729
69 Input 111100 = 60
S3=1 S4=1 S5=1 IC 8 Active
Output I60=1, verified
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
