CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1570 1 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
63
13 Logic Switch~
5 58 1772 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89956e-315 5.37752e-315
0
13 Logic Switch~
5 63 1708 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89956e-315 5.26354e-315
0
13 Logic Switch~
5 58 1912 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 513 1226 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 377 1223 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 243 1216 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 55 1574 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89956e-315 5.40342e-315
0
13 Logic Switch~
5 60 1370 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.89956e-315 5.39824e-315
0
13 Logic Switch~
5 61 1431 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.89956e-315 5.34643e-315
0
13 Logic Switch~
5 61 1027 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.89956e-315 5.37752e-315
0
13 Logic Switch~
5 60 966 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.89956e-315 5.26354e-315
0
13 Logic Switch~
5 55 1170 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 55 824 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 60 620 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 61 681 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 364 84 0 1 11
0 41
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D3
-4 -27 10 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 412 103 0 1 11
0 42
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 D2
-4 -28 10 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 463 117 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 D1
-4 -27 10 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9323 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 511 136 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 D0
-4 -27 10 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
317 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 95 377 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 MR
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3108 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 214 423 0 1 11
0 46
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 DSL
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4299 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 229 62 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 DSR
-8 -27 13 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9672 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 79 140 0 1 11
0 48
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
5.89956e-315 0
0
13 Logic Switch~
5 78 184 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
5.89956e-315 0
0
5 4013~
219 211 1808 0 6 22
0 7 2 8 6 50 5
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U9B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 8 0
1 U
9172 0 0
2
5.89956e-315 5.40342e-315
0
5 4013~
219 333 1809 0 6 22
0 7 5 8 6 51 4
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U9A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 8 0
1 U
7100 0 0
2
5.89956e-315 5.39824e-315
0
5 4013~
219 462 1808 0 6 22
0 7 4 8 6 52 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 7 0
1 U
3820 0 0
2
5.89956e-315 5.39306e-315
0
5 4013~
219 600 1808 0 6 22
0 7 3 8 6 53 2
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 7 0
1 U
7678 0 0
2
5.89956e-315 5.38788e-315
0
7 Pulser~
4 56 1845 0 10 12
0 8 54 8 55 0 0 5 5 4
7
0
0 0 4656 0
0
3 V19
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
961 0 0
2
5.89956e-315 5.36716e-315
0
14 Logic Display~
6 217 1657 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89956e-315 5.3568e-315
0
14 Logic Display~
6 339 1650 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.89956e-315 5.34643e-315
0
14 Logic Display~
6 469 1642 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.89956e-315 5.32571e-315
0
14 Logic Display~
6 687 1722 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.89956e-315 5.30499e-315
0
14 Logic Display~
6 684 1384 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.89956e-315 5.39306e-315
0
14 Logic Display~
6 466 1304 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
5.89956e-315 5.38788e-315
0
14 Logic Display~
6 336 1312 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
5.89956e-315 5.37752e-315
0
14 Logic Display~
6 214 1319 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.89956e-315 5.36716e-315
0
7 Pulser~
4 53 1507 0 10 12
0 19 56 19 57 0 0 5 5 4
7
0
0 0 4656 0
0
3 V11
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9968 0 0
2
5.89956e-315 5.3568e-315
0
5 4013~
219 597 1470 0 6 22
0 17 12 19 16 58 15
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 6 0
1 U
9281 0 0
2
5.89956e-315 5.32571e-315
0
5 4013~
219 459 1470 0 6 22
0 17 13 19 16 59 12
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 6 0
1 U
8464 0 0
2
5.89956e-315 5.30499e-315
0
5 4013~
219 330 1471 0 6 22
0 17 14 19 16 60 13
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
7168 0 0
2
5.89956e-315 5.26354e-315
0
5 4013~
219 208 1470 0 6 22
0 17 18 19 16 61 14
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 5 0
1 U
3171 0 0
2
5.89956e-315 0
0
5 4013~
219 208 1066 0 6 22
0 25 26 27 24 62 20
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 4 0
1 U
4139 0 0
2
5.89956e-315 5.26354e-315
0
5 4013~
219 330 1067 0 6 22
0 25 11 27 24 63 21
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 4 0
1 U
6435 0 0
2
5.89956e-315 0
0
5 4013~
219 459 1066 0 6 22
0 25 10 27 24 64 22
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U4B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
5283 0 0
2
5.89956e-315 5.39306e-315
0
5 4013~
219 597 1066 0 6 22
0 25 9 27 24 65 23
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U4A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
6874 0 0
2
5.89956e-315 5.38788e-315
0
7 Pulser~
4 53 1103 0 10 12
0 27 66 27 67 0 0 5 5 4
7
0
0 0 4656 0
0
2 V8
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5305 0 0
2
5.89956e-315 5.36716e-315
0
14 Logic Display~
6 214 915 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.89956e-315 5.3568e-315
0
14 Logic Display~
6 336 908 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.89956e-315 5.34643e-315
0
14 Logic Display~
6 466 900 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.89956e-315 5.32571e-315
0
14 Logic Display~
6 684 980 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.89956e-315 5.30499e-315
0
14 Logic Display~
6 684 634 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
5.89956e-315 0
0
7 Pulser~
4 53 757 0 10 12
0 35 68 35 69 0 0 5 5 4
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6118 0 0
2
5.89956e-315 0
0
5 4013~
219 597 720 0 6 22
0 30 31 35 29 70 28
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 2 0
1 U
34 0 0
2
5.89956e-315 0
0
5 4013~
219 459 720 0 6 22
0 30 32 35 29 71 31
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U3A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 2 0
1 U
6357 0 0
2
5.89956e-315 0
0
5 4013~
219 330 721 0 6 22
0 30 33 35 29 72 32
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 1 0
1 U
319 0 0
2
5.89956e-315 0
0
5 4013~
219 208 720 0 6 22
0 30 34 35 29 73 33
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 1 0
1 U
3976 0 0
2
5.89956e-315 0
0
14 Logic Display~
6 694 257 0 1 2
10 40
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
5.89956e-315 0
0
14 Logic Display~
6 655 270 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
5.89956e-315 0
0
14 Logic Display~
6 616 280 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
5.89956e-315 0
0
14 Logic Display~
6 580 288 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
5.89956e-315 0
0
7 74LS194
49 321 269 0 14 29
0 36 48 49 47 46 45 41 42 43
44 40 39 38 37
0
0 0 4848 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
842 0 0
2
5.89956e-315 0
0
7 Pulser~
4 102 242 0 10 12
0 36 74 36 75 0 0 5 5 4
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3277 0 0
2
5.89956e-315 0
0
97
1 0 2 0 0 4224 0 33 0 0 17 3
687 1740
122 1740
122 1772
0 2 3 0 0 4096 0 0 28 7 0 2
514 1772
576 1772
0 2 4 0 0 8192 0 0 27 6 0 3
387 1773
387 1772
438 1772
0 2 5 0 0 8192 0 0 26 5 0 3
276 1772
276 1773
309 1773
6 1 5 0 0 8320 0 25 30 0 0 4
235 1772
276 1772
276 1675
217 1675
6 1 4 0 0 8320 0 26 31 0 0 4
357 1773
387 1773
387 1668
339 1668
6 1 3 0 0 8320 0 27 32 0 0 4
486 1772
514 1772
514 1660
469 1660
6 1 2 0 0 0 0 28 33 0 0 3
624 1772
687 1772
687 1740
0 4 6 0 0 4096 0 0 28 10 0 3
462 1912
600 1912
600 1814
0 4 6 0 0 0 0 0 27 11 0 3
333 1912
462 1912
462 1814
0 4 6 0 0 0 0 0 26 12 0 3
211 1912
333 1912
333 1815
1 4 6 0 0 4224 0 3 25 0 0 3
70 1912
211 1912
211 1814
0 1 7 0 0 4224 0 0 28 14 0 3
462 1708
600 1708
600 1751
0 1 7 0 0 0 0 0 27 15 0 3
333 1708
462 1708
462 1751
0 1 7 0 0 0 0 0 26 16 0 3
211 1708
333 1708
333 1752
1 1 7 0 0 0 0 2 25 0 0 3
75 1708
211 1708
211 1751
1 2 2 0 0 0 0 1 25 0 0 2
70 1772
187 1772
0 3 8 0 0 4224 0 0 28 19 0 3
438 1836
576 1836
576 1790
0 3 8 0 0 0 0 0 27 20 0 3
309 1836
438 1836
438 1790
0 3 8 0 0 0 0 0 26 22 0 3
187 1836
309 1836
309 1791
1 0 8 0 0 0 0 29 0 0 22 5
32 1836
23 1836
23 1811
118 1811
118 1836
3 3 8 0 0 0 0 29 25 0 0 3
80 1836
187 1836
187 1790
1 2 9 0 0 8320 0 4 46 0 0 4
525 1226
565 1226
565 1030
573 1030
1 2 10 0 0 8320 0 5 45 0 0 4
389 1223
423 1223
423 1030
435 1030
1 2 11 0 0 8320 0 6 44 0 0 4
255 1216
288 1216
288 1031
306 1031
0 2 12 0 0 4096 0 0 39 31 0 2
511 1434
573 1434
0 2 13 0 0 8192 0 0 40 30 0 3
384 1435
384 1434
435 1434
0 2 14 0 0 8192 0 0 41 29 0 3
273 1434
273 1435
306 1435
6 1 14 0 0 8320 0 42 37 0 0 4
232 1434
273 1434
273 1337
214 1337
6 1 13 0 0 8320 0 41 36 0 0 4
354 1435
384 1435
384 1330
336 1330
6 1 12 0 0 8320 0 40 35 0 0 4
483 1434
511 1434
511 1322
466 1322
6 1 15 0 0 4224 0 39 34 0 0 3
621 1434
684 1434
684 1402
0 4 16 0 0 4096 0 0 39 34 0 3
459 1574
597 1574
597 1476
0 4 16 0 0 0 0 0 40 35 0 3
330 1574
459 1574
459 1476
0 4 16 0 0 0 0 0 41 36 0 3
208 1574
330 1574
330 1477
1 4 16 0 0 4224 0 7 42 0 0 3
67 1574
208 1574
208 1476
0 1 17 0 0 4224 0 0 39 38 0 3
459 1370
597 1370
597 1413
0 1 17 0 0 0 0 0 40 39 0 3
330 1370
459 1370
459 1413
0 1 17 0 0 0 0 0 41 40 0 3
208 1370
330 1370
330 1414
1 1 17 0 0 0 0 8 42 0 0 3
72 1370
208 1370
208 1413
1 2 18 0 0 8320 0 9 42 0 0 3
73 1431
73 1434
184 1434
0 3 19 0 0 4224 0 0 39 43 0 3
435 1498
573 1498
573 1452
0 3 19 0 0 0 0 0 40 44 0 3
306 1498
435 1498
435 1452
0 3 19 0 0 0 0 0 41 46 0 3
184 1498
306 1498
306 1453
1 0 19 0 0 0 0 38 0 0 46 5
29 1498
20 1498
20 1473
115 1473
115 1498
3 3 19 0 0 0 0 38 42 0 0 3
77 1498
184 1498
184 1452
6 1 20 0 0 8320 0 43 48 0 0 4
232 1030
273 1030
273 933
214 933
6 1 21 0 0 8320 0 44 49 0 0 4
354 1031
384 1031
384 926
336 926
6 1 22 0 0 8320 0 45 50 0 0 4
483 1030
511 1030
511 918
466 918
6 1 23 0 0 4224 0 46 51 0 0 3
621 1030
684 1030
684 998
0 4 24 0 0 4096 0 0 46 52 0 3
459 1170
597 1170
597 1072
0 4 24 0 0 0 0 0 45 53 0 3
330 1170
459 1170
459 1072
0 4 24 0 0 0 0 0 44 54 0 3
208 1170
330 1170
330 1073
1 4 24 0 0 4224 0 12 43 0 0 3
67 1170
208 1170
208 1072
0 1 25 0 0 4224 0 0 46 56 0 3
459 966
597 966
597 1009
0 1 25 0 0 0 0 0 45 57 0 3
330 966
459 966
459 1009
0 1 25 0 0 0 0 0 44 58 0 3
208 966
330 966
330 1010
1 1 25 0 0 0 0 11 43 0 0 3
72 966
208 966
208 1009
1 2 26 0 0 8320 0 10 43 0 0 3
73 1027
73 1030
184 1030
0 3 27 0 0 4224 0 0 46 61 0 3
435 1094
573 1094
573 1048
0 3 27 0 0 0 0 0 45 62 0 3
306 1094
435 1094
435 1048
0 3 27 0 0 0 0 0 44 64 0 3
184 1094
306 1094
306 1049
1 0 27 0 0 0 0 47 0 0 64 5
29 1094
20 1094
20 1069
115 1069
115 1094
3 3 27 0 0 0 0 47 43 0 0 3
77 1094
184 1094
184 1048
6 1 28 0 0 4224 0 54 52 0 0 3
621 684
684 684
684 652
0 4 29 0 0 4096 0 0 54 67 0 3
459 824
597 824
597 726
0 4 29 0 0 0 0 0 55 68 0 3
330 824
459 824
459 726
0 4 29 0 0 0 0 0 56 69 0 3
208 824
330 824
330 727
1 4 29 0 0 4224 0 13 57 0 0 3
67 824
208 824
208 726
0 1 30 0 0 4224 0 0 54 71 0 3
459 620
597 620
597 663
0 1 30 0 0 0 0 0 55 72 0 3
330 620
459 620
459 663
0 1 30 0 0 0 0 0 56 73 0 3
208 620
330 620
330 664
1 1 30 0 0 0 0 14 57 0 0 3
72 620
208 620
208 663
6 2 31 0 0 4224 0 55 54 0 0 2
483 684
573 684
6 2 32 0 0 8320 0 56 55 0 0 3
354 685
354 684
435 684
6 2 33 0 0 8320 0 57 56 0 0 3
232 684
232 685
306 685
1 2 34 0 0 8320 0 15 57 0 0 3
73 681
73 684
184 684
0 3 35 0 0 4224 0 0 54 79 0 3
435 748
573 748
573 702
0 3 35 0 0 0 0 0 55 80 0 3
306 748
435 748
435 702
0 3 35 0 0 0 0 0 56 82 0 3
184 748
306 748
306 703
1 0 35 0 0 0 0 53 0 0 82 5
29 748
20 748
20 723
115 723
115 748
3 3 35 0 0 0 0 53 57 0 0 3
77 748
184 748
184 702
3 0 36 0 0 4096 0 63 0 0 84 2
126 233
153 233
1 1 36 0 0 16512 0 63 62 0 0 5
78 233
78 200
153 200
153 233
289 233
1 14 37 0 0 8320 0 61 62 0 0 3
580 306
580 305
353 305
1 13 38 0 0 8320 0 60 62 0 0 3
616 298
616 296
353 296
1 12 39 0 0 8320 0 59 62 0 0 3
655 288
655 287
353 287
1 11 40 0 0 8320 0 58 62 0 0 3
694 275
694 278
353 278
1 7 41 0 0 4224 0 16 62 0 0 3
376 84
376 233
353 233
1 8 42 0 0 4224 0 17 62 0 0 3
424 103
424 242
353 242
1 9 43 0 0 4224 0 18 62 0 0 3
475 117
475 251
353 251
1 10 44 0 0 8320 0 19 62 0 0 3
523 136
523 260
353 260
1 6 45 0 0 4224 0 20 62 0 0 4
107 377
261 377
261 305
283 305
1 5 46 0 0 4224 0 21 62 0 0 3
226 423
226 287
289 287
1 4 47 0 0 4224 0 22 62 0 0 3
241 62
241 278
289 278
1 2 48 0 0 4224 0 23 62 0 0 4
91 140
231 140
231 251
289 251
1 3 49 0 0 4224 0 24 62 0 0 4
90 184
219 184
219 260
289 260
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
