CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 253 235 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44010.8 10
0
13 Logic Switch~
5 266 171 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
44010.8 9
0
13 Logic Switch~
5 264 134 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44010.8 8
0
13 Logic Switch~
5 259 88 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44010.8 7
0
13 Logic Switch~
5 259 50 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44010.8 6
0
13 Logic Switch~
5 45 121 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-4 -28 3 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
44010.8 8
0
13 Logic Switch~
5 47 180 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44010.8 7
0
13 Logic Switch~
5 29 219 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -25 4 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44010.8 2
0
13 Logic Switch~
5 36 255 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
44010.8 1
0
13 Logic Switch~
5 46 94 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
5.89944e-315 0
0
13 Logic Switch~
5 44 39 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
5.89944e-315 0
0
14 Logic Display~
6 364 218 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
44010.8 5
0
9 Inverter~
13 308 236 0 2 22
0 2 3
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
3536 0 0
2
44010.8 4
0
14 Logic Display~
6 405 129 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44010.8 3
0
14 Logic Display~
6 400 42 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
44010.8 2
0
9 2-In XOR~
219 342 147 0 3 22
0 5 4 6
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3670 0 0
2
44010.8 1
0
9 2-In NOR~
219 321 63 0 3 22
0 9 8 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 NOR
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
5616 0 0
2
44010.8 0
0
8 2-In OR~
219 110 153 0 3 22
0 13 14 15
0
0 0 624 0
5 74F32
-18 -24 17 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
44010.8 18
0
14 Logic Display~
6 181 135 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
44010.8 17
0
10 2-In NAND~
219 127 224 0 3 22
0 11 10 12
0
0 0 624 0
4 7400
-7 -24 21 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3108 0 0
2
44010.8 16
0
14 Logic Display~
6 188 206 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
44010.8 13
0
14 Logic Display~
6 175 50 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89944e-315 0
0
9 2-In AND~
219 118 68 0 3 22
0 17 16 18
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7876 0 0
2
5.89944e-315 0
0
17
1 1 2 0 0 8336 0 13 1 0 0 3
293 236
293 235
265 235
1 2 3 0 0 4240 0 12 13 0 0 2
364 236
329 236
2 1 4 0 0 4240 0 16 2 0 0 3
326 156
278 156
278 171
1 1 5 0 0 4240 0 16 3 0 0 3
326 138
276 138
276 134
1 3 6 0 0 4240 0 14 16 0 0 2
405 147
375 147
1 3 7 0 0 8336 0 15 17 0 0 3
400 60
400 63
360 63
2 1 8 0 0 4240 0 17 4 0 0 3
308 72
271 72
271 88
1 1 9 0 0 4240 0 17 5 0 0 3
308 54
271 54
271 50
2 1 10 0 0 4224 0 20 9 0 0 3
103 233
48 233
48 255
1 1 11 0 0 4224 0 20 8 0 0 3
103 215
41 215
41 219
1 3 12 0 0 4224 0 21 20 0 0 2
188 224
154 224
1 1 13 0 0 4224 0 18 6 0 0 4
97 144
58 144
58 121
57 121
2 1 14 0 0 4224 0 18 7 0 0 3
97 162
59 162
59 180
1 3 15 0 0 4224 0 19 18 0 0 2
181 153
143 153
1 2 16 0 0 4224 0 10 23 0 0 4
58 94
79 94
79 77
94 77
1 1 17 0 0 4224 0 11 23 0 0 4
56 39
79 39
79 59
94 59
1 3 18 0 0 4224 0 22 23 0 0 2
175 68
139 68
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
315 163 330 187
318 165 326 181
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
278 212 293 236
281 214 289 230
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
303 31 318 55
306 33 314 49
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
303 79 318 103
306 81 314 97
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
311 111 332 132
317 117 325 132
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
92 83 107 107
95 85 103 101
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
91 168 106 192
94 170 102 186
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
90 35 105 59
93 37 101 53
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
91 112 106 136
94 114 102 130
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
100 241 115 265
103 243 111 259
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
99 192 114 216
102 194 110 210
1 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
