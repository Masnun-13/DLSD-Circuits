CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 1 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 120 645 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 PRE3
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
659 0 0
2
5.89957e-315 5.41378e-315
0
13 Logic Switch~
5 122 767 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 CLR3
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3800 0 0
2
5.89957e-315 5.4086e-315
0
13 Logic Switch~
5 91 613 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 L9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6792 0 0
2
5.89957e-315 5.40342e-315
0
13 Logic Switch~
5 57 514 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 M
-2 -26 5 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3701 0 0
2
5.89957e-315 5.39824e-315
0
13 Logic Switch~
5 127 348 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 PRE2
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6316 0 0
2
5.89957e-315 5.30499e-315
0
13 Logic Switch~
5 93 470 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 CLR2
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8734 0 0
2
5.89957e-315 5.26354e-315
0
13 Logic Switch~
5 62 319 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 L8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7988 0 0
2
5.89957e-315 0
0
13 Logic Switch~
5 89 77 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 L1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3217 0 0
2
5.89957e-315 5.39306e-315
0
13 Logic Switch~
5 120 231 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 CLR1
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3965 0 0
2
5.89957e-315 5.37752e-315
0
13 Logic Switch~
5 118 109 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 PRE1
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8239 0 0
2
5.89957e-315 5.36716e-315
0
9 2-In XOR~
219 501 743 0 3 22
0 7 5 4
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
828 0 0
2
5.89957e-315 5.39306e-315
0
9 2-In AND~
219 569 673 0 3 22
0 3 4 2
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
6187 0 0
2
5.89957e-315 5.38788e-315
0
9 2-In XOR~
219 317 673 0 3 22
0 7 6 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
7107 0 0
2
5.89957e-315 5.37752e-315
0
5 4027~
219 630 709 0 7 32
0 9 2 8 2 10 31 11
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
6433 0 0
2
5.89957e-315 5.36716e-315
0
5 4027~
219 436 709 0 7 32
0 9 3 8 3 10 32 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8559 0 0
2
5.89957e-315 5.3568e-315
0
5 4027~
219 225 709 0 7 32
0 9 12 8 12 10 33 6
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3674 0 0
2
5.89957e-315 5.34643e-315
0
14 Logic Display~
6 722 585 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5697 0 0
2
5.89957e-315 5.32571e-315
0
14 Logic Display~
6 501 588 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3805 0 0
2
5.89957e-315 5.30499e-315
0
14 Logic Display~
6 286 590 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5219 0 0
2
5.89957e-315 5.26354e-315
0
7 Pulser~
4 89 691 0 10 12
0 34 8 35 8 0 0 5 5 3
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3795 0 0
2
5.89957e-315 0
0
5 4027~
219 601 415 0 7 32
0 17 13 16 13 18 36 19
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U3B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
3637 0 0
2
5.89957e-315 5.43192e-315
0
5 4027~
219 407 415 0 7 32
0 17 14 16 14 18 15 20
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U4A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 4 0
1 U
3226 0 0
2
5.89957e-315 5.42933e-315
0
5 4027~
219 196 415 0 7 32
0 17 22 16 22 18 14 21
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U4B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 4 0
1 U
6966 0 0
2
5.89957e-315 5.42414e-315
0
14 Logic Display~
6 287 286 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9796 0 0
2
5.89957e-315 5.41896e-315
0
7 Pulser~
4 60 397 0 10 12
0 16 37 16 38 0 0 5 5 3
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5952 0 0
2
5.89957e-315 5.41378e-315
0
14 Logic Display~
6 473 291 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3649 0 0
2
5.89957e-315 5.4086e-315
0
14 Logic Display~
6 694 289 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3716 0 0
2
5.89957e-315 5.40342e-315
0
9 2-In AND~
219 528 379 0 3 22
0 15 14 13
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4797 0 0
2
5.89957e-315 5.39824e-315
0
9 2-In AND~
219 538 137 0 3 22
0 25 24 23
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
4681 0 0
2
5.89957e-315 0
0
7 Pulser~
4 87 155 0 10 12
0 39 26 40 26 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9730 0 0
2
5.89957e-315 5.47077e-315
0
14 Logic Display~
6 284 54 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9874 0 0
2
5.89957e-315 5.46818e-315
0
14 Logic Display~
6 499 52 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
364 0 0
2
5.89957e-315 5.46559e-315
0
14 Logic Display~
6 720 49 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3656 0 0
2
5.89957e-315 5.463e-315
0
5 4027~
219 223 173 0 7 32
0 27 30 26 30 28 41 25
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U6A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 6 0
1 U
3131 0 0
2
5.89957e-315 5.45005e-315
0
5 4027~
219 434 173 0 7 32
0 27 25 26 25 28 42 24
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
6772 0 0
2
5.89957e-315 5.44746e-315
0
5 4027~
219 628 173 0 7 32
0 27 23 26 23 28 43 29
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
9557 0 0
2
5.89957e-315 5.44487e-315
0
67
0 4 2 0 0 4224 0 0 14 2 0 3
600 673
600 691
606 691
3 2 2 0 0 128 0 12 14 0 0 2
590 673
606 673
0 1 3 0 0 8320 0 0 12 5 0 3
383 673
383 664
545 664
0 4 3 0 0 0 0 0 15 5 0 3
399 673
399 691
412 691
3 2 3 0 0 0 0 13 15 0 0 2
350 673
412 673
3 2 4 0 0 8320 0 11 12 0 0 3
534 743
545 743
545 682
0 2 5 0 0 4224 0 0 11 22 0 3
472 673
472 752
485 752
0 2 6 0 0 8192 0 0 13 23 0 3
274 673
274 682
301 682
1 0 7 0 0 8320 0 11 0 0 10 4
485 734
361 734
361 514
274 514
1 1 7 0 0 0 0 4 13 0 0 4
69 514
274 514
274 664
301 664
3 0 8 0 0 8192 0 15 0 0 12 3
412 682
380 682
380 722
0 3 8 0 0 8320 0 0 14 14 0 5
165 682
165 722
589 722
589 682
606 682
0 4 8 0 0 0 0 0 20 14 0 3
133 682
133 691
119 691
2 3 8 0 0 0 0 20 16 0 0 6
59 691
50 691
50 658
133 658
133 682
201 682
0 1 9 0 0 4096 0 0 14 16 0 3
436 645
630 645
630 652
0 1 9 0 0 4224 0 0 15 17 0 3
225 645
436 645
436 652
1 1 9 0 0 0 0 1 16 0 0 3
132 645
225 645
225 652
0 5 10 0 0 4096 0 0 14 19 0 3
436 767
630 767
630 715
0 5 10 0 0 4224 0 0 15 20 0 3
225 767
436 767
436 715
1 5 10 0 0 0 0 2 16 0 0 3
134 767
225 767
225 715
7 1 11 0 0 8320 0 14 17 0 0 3
654 673
722 673
722 603
7 1 5 0 0 0 0 15 18 0 0 3
460 673
501 673
501 606
7 1 6 0 0 8320 0 16 19 0 0 3
249 673
286 673
286 608
0 4 12 0 0 4096 0 0 16 25 0 3
192 672
192 691
201 691
1 2 12 0 0 4224 0 3 16 0 0 4
103 613
192 613
192 673
201 673
0 4 13 0 0 4096 0 0 21 27 0 3
566 379
566 397
577 397
3 2 13 0 0 4224 0 28 21 0 0 2
549 379
577 379
0 2 14 0 0 8320 0 0 28 31 0 5
314 397
314 419
500 419
500 388
504 388
6 1 15 0 0 4224 0 22 28 0 0 4
437 397
486 397
486 370
504 370
0 2 14 0 0 0 0 0 22 31 0 3
349 397
349 379
383 379
6 4 14 0 0 0 0 23 22 0 0 2
226 397
383 397
3 0 16 0 0 8192 0 22 0 0 33 3
383 388
363 388
363 427
0 3 16 0 0 8320 0 0 21 46 0 5
136 388
136 427
557 427
557 388
577 388
0 1 17 0 0 8192 0 0 23 36 0 3
195 348
196 348
196 358
0 1 17 0 0 0 0 0 22 36 0 2
407 348
407 358
1 1 17 0 0 4224 0 5 21 0 0 3
139 348
601 348
601 358
0 5 18 0 0 4096 0 0 21 38 0 3
407 470
601 470
601 421
0 5 18 0 0 4224 0 0 22 39 0 3
196 470
407 470
407 421
1 5 18 0 0 0 0 6 23 0 0 3
105 470
196 470
196 421
7 1 19 0 0 8320 0 21 27 0 0 3
625 379
694 379
694 307
7 1 20 0 0 8320 0 22 26 0 0 3
431 379
473 379
473 309
7 1 21 0 0 8320 0 23 24 0 0 3
220 379
287 379
287 304
0 4 22 0 0 4096 0 0 23 44 0 3
163 378
163 397
172 397
1 2 22 0 0 4224 0 7 23 0 0 4
74 319
163 319
163 379
172 379
1 0 16 0 0 0 0 25 0 0 46 5
36 388
27 388
27 362
98 362
98 388
3 3 16 0 0 0 0 25 23 0 0 2
84 388
172 388
0 4 23 0 0 4096 0 0 36 48 0 3
591 137
591 155
604 155
3 2 23 0 0 4224 0 29 36 0 0 2
559 137
604 137
0 2 24 0 0 8192 0 0 29 64 0 3
485 137
485 146
514 146
1 0 25 0 0 4224 0 29 0 0 65 2
514 128
284 128
3 0 26 0 0 8192 0 35 0 0 52 3
410 146
371 146
371 186
0 3 26 0 0 8320 0 0 36 56 0 5
164 146
164 186
558 186
558 146
604 146
0 4 25 0 0 0 0 0 35 54 0 3
400 137
400 155
410 155
0 2 25 0 0 0 0 0 35 65 0 2
282 137
410 137
0 4 26 0 0 0 0 0 30 56 0 3
131 146
131 155
117 155
2 3 26 0 0 0 0 30 34 0 0 6
57 155
48 155
48 122
131 122
131 146
199 146
0 1 27 0 0 4096 0 0 36 58 0 3
434 109
628 109
628 116
0 1 27 0 0 4224 0 0 35 59 0 3
223 109
434 109
434 116
1 1 27 0 0 0 0 10 34 0 0 3
130 109
223 109
223 116
0 5 28 0 0 4096 0 0 36 61 0 3
434 231
628 231
628 179
0 5 28 0 0 4224 0 0 35 62 0 3
223 231
434 231
434 179
1 5 28 0 0 0 0 9 34 0 0 3
132 231
223 231
223 179
7 1 29 0 0 8320 0 36 33 0 0 3
652 137
720 137
720 67
7 1 24 0 0 8320 0 35 32 0 0 3
458 137
499 137
499 70
7 1 25 0 0 0 0 34 31 0 0 3
247 137
284 137
284 72
0 4 30 0 0 4096 0 0 34 67 0 3
190 136
190 155
199 155
1 2 30 0 0 4224 0 8 34 0 0 4
101 77
190 77
190 137
199 137
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
