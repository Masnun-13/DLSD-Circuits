CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 110 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 488 348 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44074 0
0
13 Logic Switch~
5 451 418 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44074 1
0
13 Logic Switch~
5 834 230 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
44074 2
0
13 Logic Switch~
5 528 121 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
44074 3
0
13 Logic Switch~
5 514 237 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
44074 4
0
13 Logic Switch~
5 512 541 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
44074 5
0
13 Logic Switch~
5 526 425 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
44074 6
0
13 Logic Switch~
5 824 415 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
44074 7
0
13 Logic Switch~
5 336 414 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
44074 8
0
13 Logic Switch~
5 38 424 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
44074 9
0
13 Logic Switch~
5 24 540 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
44074 10
0
13 Logic Switch~
5 26 236 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
44074 11
0
13 Logic Switch~
5 40 120 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
44074 12
0
13 Logic Switch~
5 346 229 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
44074 13
0
7 74LS153
119 792 314 0 14 29
0 19 18 17 16 2 3 9 5 8
7 15 4 13 6
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
3835 0 0
2
44074 14
0
9 2-In AND~
219 627 305 0 3 22
0 12 14 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3670 0 0
2
44074 15
0
8 2-In OR~
219 623 228 0 3 22
0 12 14 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
5616 0 0
2
44074 16
0
9 2-In XOR~
219 628 174 0 3 22
0 12 14 18
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9323 0 0
2
44074 17
0
9 Inverter~
13 626 121 0 2 22
0 12 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
317 0 0
2
44074 18
0
14 Logic Display~
6 944 320 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44074 19
0
9 Inverter~
13 624 425 0 2 22
0 10 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
4299 0 0
2
44074 20
0
9 2-In XOR~
219 628 479 0 3 22
0 10 11 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9672 0 0
2
44074 21
0
8 2-In OR~
219 621 532 0 3 22
0 10 11 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7876 0 0
2
44074 22
0
9 2-In AND~
219 630 583 0 3 22
0 10 11 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6369 0 0
2
44074 23
0
14 Logic Display~
6 923 322 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
44074 24
0
14 Logic Display~
6 965 316 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
44074 25
0
9 2-In AND~
219 142 582 0 3 22
0 26 27 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3820 0 0
2
44074 26
0
8 2-In OR~
219 133 531 0 3 22
0 26 27 24
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7678 0 0
2
44074 27
0
9 2-In XOR~
219 140 478 0 3 22
0 26 27 21
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
961 0 0
2
44074 28
0
9 Inverter~
13 136 424 0 2 22
0 26 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3178 0 0
2
44074 29
0
14 Logic Display~
6 985 316 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
44074 30
0
9 Inverter~
13 138 120 0 2 22
0 28 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3951 0 0
2
44074 31
0
9 2-In XOR~
219 140 173 0 3 22
0 28 30 34
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8885 0 0
2
44074 32
0
8 2-In OR~
219 135 227 0 3 22
0 28 30 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3780 0 0
2
44074 33
0
9 2-In AND~
219 139 304 0 3 22
0 28 30 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9265 0 0
2
44074 34
0
7 74LS153
119 304 313 0 14 29
0 35 34 33 32 2 3 25 21 24
23 31 20 29 22
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
9442 0 0
2
44074 35
0
56
1 5 2 0 0 8320 0 1 36 0 0 5
500 348
500 384
209 384
209 313
272 313
1 6 3 0 0 12288 0 2 15 0 0 6
463 418
485 418
485 368
684 368
684 323
760 323
1 6 3 0 0 8320 0 2 36 0 0 5
463 418
463 441
236 441
236 322
272 322
1 5 2 0 0 0 0 1 15 0 0 4
500 348
655 348
655 314
760 314
1 12 4 0 0 8320 0 8 15 0 0 4
836 415
850 415
850 359
830 359
8 3 5 0 0 8320 0 15 22 0 0 4
760 341
744 341
744 479
661 479
1 14 6 0 0 8320 0 25 15 0 0 3
923 340
923 341
824 341
3 10 7 0 0 8320 0 24 15 0 0 3
651 583
760 583
760 359
3 9 8 0 0 8320 0 23 15 0 0 4
654 532
750 532
750 350
760 350
2 7 9 0 0 8320 0 21 15 0 0 4
645 425
737 425
737 332
760 332
0 1 10 0 0 4096 0 0 22 13 0 2
569 470
612 470
0 1 10 0 0 0 0 0 23 13 0 2
569 523
608 523
0 1 10 0 0 4224 0 0 24 14 0 3
569 425
569 574
606 574
1 1 10 0 0 0 0 7 21 0 0 2
538 425
609 425
1 2 11 0 0 8192 0 6 24 0 0 3
524 541
524 592
606 592
1 2 11 0 0 4096 0 6 23 0 0 2
524 541
608 541
1 2 11 0 0 8320 0 6 22 0 0 3
524 541
524 488
612 488
0 1 12 0 0 8192 0 0 18 20 0 3
571 166
571 165
612 165
0 1 12 0 0 0 0 0 17 20 0 2
571 219
610 219
0 1 12 0 0 4224 0 0 16 21 0 3
571 121
571 296
603 296
1 1 12 0 0 0 0 4 19 0 0 2
540 121
611 121
1 13 13 0 0 4224 0 20 15 0 0 4
944 338
839 338
839 296
824 296
1 2 14 0 0 4096 0 5 16 0 0 3
526 237
526 314
603 314
1 2 14 0 0 4096 0 5 17 0 0 2
526 237
610 237
1 2 14 0 0 8320 0 5 18 0 0 3
526 237
526 183
612 183
1 11 15 0 0 4224 0 3 15 0 0 3
846 230
846 278
830 278
3 4 16 0 0 4224 0 16 15 0 0 2
648 305
760 305
3 3 17 0 0 12416 0 17 15 0 0 4
656 228
659 228
659 296
760 296
3 2 18 0 0 8320 0 18 15 0 0 4
661 174
668 174
668 287
760 287
2 1 19 0 0 8320 0 19 15 0 0 4
647 121
691 121
691 278
760 278
1 12 20 0 0 8320 0 9 36 0 0 4
348 414
362 414
362 358
342 358
8 3 21 0 0 8320 0 36 29 0 0 4
272 340
256 340
256 478
173 478
1 14 22 0 0 8320 0 26 36 0 0 3
965 334
965 340
336 340
3 10 23 0 0 8320 0 27 36 0 0 3
163 582
272 582
272 358
3 9 24 0 0 8320 0 28 36 0 0 4
166 531
262 531
262 349
272 349
2 7 25 0 0 8320 0 30 36 0 0 4
157 424
249 424
249 331
272 331
0 1 26 0 0 4096 0 0 29 39 0 2
81 469
124 469
0 1 26 0 0 0 0 0 28 39 0 2
81 522
120 522
0 1 26 0 0 4224 0 0 27 40 0 3
81 424
81 573
118 573
1 1 26 0 0 0 0 10 30 0 0 2
50 424
121 424
1 2 27 0 0 8192 0 11 27 0 0 3
36 540
36 591
118 591
1 2 27 0 0 4096 0 11 28 0 0 2
36 540
120 540
1 2 27 0 0 8320 0 11 29 0 0 3
36 540
36 487
124 487
0 1 28 0 0 8192 0 0 33 46 0 3
83 165
83 164
124 164
0 1 28 0 0 0 0 0 34 46 0 2
83 218
122 218
0 1 28 0 0 4224 0 0 35 47 0 3
83 120
83 295
115 295
1 1 28 0 0 0 0 13 32 0 0 2
52 120
123 120
1 13 29 0 0 4224 0 31 36 0 0 4
985 334
351 334
351 295
336 295
1 2 30 0 0 4096 0 12 35 0 0 3
38 236
38 313
115 313
1 2 30 0 0 4096 0 12 34 0 0 2
38 236
122 236
1 2 30 0 0 8320 0 12 33 0 0 3
38 236
38 182
124 182
1 11 31 0 0 4224 0 14 36 0 0 3
358 229
358 277
342 277
3 4 32 0 0 4224 0 35 36 0 0 2
160 304
272 304
3 3 33 0 0 12416 0 34 36 0 0 4
168 227
171 227
171 295
272 295
3 2 34 0 0 8320 0 33 36 0 0 4
173 173
180 173
180 286
272 286
2 1 35 0 0 8320 0 32 36 0 0 4
159 120
203 120
203 277
272 277
44
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
106 91 133 113
115 99 123 115
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
109 134 136 156
118 142 126 158
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
105 189 132 211
114 197 122 213
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
104 265 131 287
113 273 121 289
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
104 316 127 338
111 324 119 340
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
108 239 131 261
115 247 123 263
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
114 177 137 199
121 185 129 201
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
153 95 176 117
160 103 168 119
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
102 398 127 420
110 405 118 421
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
157 308 182 330
165 315 173 331
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
157 205 182 227
165 212 173 228
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
166 151 191 173
174 158 182 174
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
147 397 172 419
155 405 163 421
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
107 444 132 466
115 452 123 468
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
111 493 136 515
119 501 127 517
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
105 551 130 573
113 559 121 575
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
106 482 131 504
114 489 122 505
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
107 536 132 558
115 544 123 560
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
106 591 131 613
114 598 122 614
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
593 93 618 115
601 100 609 116
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
639 97 662 119
646 105 654 121
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
164 453 187 475
171 461 179 477
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
158 505 181 527
165 513 173 529
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
154 560 177 582
161 568 169 584
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
585 139 618 161
593 146 609 162
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
584 196 617 218
592 203 608 219
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
585 274 618 296
593 281 609 297
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
588 177 615 199
597 185 605 201
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
590 236 617 258
599 244 607 260
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
588 309 615 331
597 317 605 333
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
591 397 618 419
600 405 608 421
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
635 399 660 421
643 406 651 422
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
638 286 663 308
646 293 654 309
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
641 205 666 227
649 212 657 228
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
648 150 673 172
656 157 664 173
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
587 444 622 466
596 451 612 467
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
582 497 617 519
591 504 607 520
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
581 550 616 572
590 557 606 573
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
591 481 626 503
600 488 616 504
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
586 536 621 558
595 543 611 559
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
587 594 622 616
596 601 612 617
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
640 558 675 580
649 565 665 581
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
645 506 680 528
654 513 670 529
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
652 451 687 473
661 458 677 474
2 11
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
