CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 50 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
142
13 Logic Switch~
5 33 411 0 1 11
0 67
0
0 0 21360 0
2 0V
-6 -17 8 -9
1 E
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44105.3 0
0
13 Logic Switch~
5 32 367 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
1 D
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44105.3 0
0
13 Logic Switch~
5 67 163 0 1 11
0 132
0
0 0 21360 0
2 0V
-9 -15 5 -7
1 C
-4 -29 3 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44105.3 0
0
13 Logic Switch~
5 66 214 0 10 11
0 131 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
44105.3 0
0
13 Logic Switch~
5 63 263 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -17 8 -9
1 A
-3 -28 4 -20
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
44105.3 0
0
9 Inverter~
13 1646 542 0 2 22
0 2 3
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
5572 0 0
2
44105.3 41
0
14 Logic Display~
6 1649 508 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out32
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
44105.3 40
0
9 Inverter~
13 1599 541 0 2 22
0 4 5
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
7361 0 0
2
44105.3 39
0
14 Logic Display~
6 1602 507 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out33
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
44105.3 38
0
9 Inverter~
13 1554 542 0 2 22
0 6 7
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 6 0
1 U
972 0 0
2
44105.3 37
0
14 Logic Display~
6 1557 508 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out34
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
44105.3 36
0
9 Inverter~
13 1504 544 0 2 22
0 8 9
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
9998 0 0
2
44105.3 35
0
14 Logic Display~
6 1507 510 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out35
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
44105.3 34
0
9 Inverter~
13 1450 541 0 2 22
0 10 11
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
4597 0 0
2
44105.3 33
0
14 Logic Display~
6 1453 507 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out36
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
44105.3 32
0
9 Inverter~
13 1404 542 0 2 22
0 12 13
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
3670 0 0
2
44105.3 31
0
14 Logic Display~
6 1407 508 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out37
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
44105.3 30
0
9 Inverter~
13 1355 541 0 2 22
0 14 15
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 7 0
1 U
9323 0 0
2
44105.3 29
0
14 Logic Display~
6 1358 507 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out38
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
44105.3 28
0
9 Inverter~
13 1312 539 0 2 22
0 16 17
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 7 0
1 U
3108 0 0
2
44105.3 27
0
14 Logic Display~
6 1315 505 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out39
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
44105.3 26
0
9 Inverter~
13 1646 405 0 2 22
0 18 19
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 7 0
1 U
9672 0 0
2
44105.3 25
0
14 Logic Display~
6 1649 371 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out40
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
44105.3 24
0
9 Inverter~
13 1599 404 0 2 22
0 20 21
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
6369 0 0
2
44105.3 23
0
14 Logic Display~
6 1602 370 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out41
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9172 0 0
2
44105.3 22
0
9 Inverter~
13 1556 403 0 2 22
0 22 23
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
7100 0 0
2
44105.3 21
0
14 Logic Display~
6 1559 369 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out42
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3820 0 0
2
44105.3 20
0
9 Inverter~
13 1505 405 0 2 22
0 24 25
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
7678 0 0
2
44105.3 19
0
14 Logic Display~
6 1508 371 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out43
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
961 0 0
2
44105.3 18
0
9 Inverter~
13 1451 406 0 2 22
0 26 27
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
3178 0 0
2
44105.3 17
0
14 Logic Display~
6 1454 372 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out44
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
44105.3 16
0
9 Inverter~
13 1405 405 0 2 22
0 28 29
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3951 0 0
2
44105.3 15
0
14 Logic Display~
6 1408 371 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out45
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
44105.3 14
0
9 Inverter~
13 1356 405 0 2 22
0 30 31
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U12F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3780 0 0
2
44105.3 13
0
14 Logic Display~
6 1359 371 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out46
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
44105.3 12
0
9 Inverter~
13 1313 406 0 2 22
0 32 33
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
9442 0 0
2
44105.3 11
0
14 Logic Display~
6 1316 372 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out47
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9424 0 0
2
44105.3 10
0
9 Inverter~
13 1642 269 0 2 22
0 34 35
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
9968 0 0
2
44105.3 9
0
14 Logic Display~
6 1645 235 0 1 2
10 35
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out48
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9281 0 0
2
44105.3 8
0
9 Inverter~
13 1595 267 0 2 22
0 36 37
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
8464 0 0
2
44105.3 7
0
14 Logic Display~
6 1598 233 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out49
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
44105.3 6
0
9 Inverter~
13 1552 267 0 2 22
0 38 39
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
3171 0 0
2
44105.3 5
0
14 Logic Display~
6 1555 233 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out50
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4139 0 0
2
44105.3 4
0
9 Inverter~
13 1501 268 0 2 22
0 40 41
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
6435 0 0
2
44105.3 3
0
14 Logic Display~
6 1504 234 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out51
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5283 0 0
2
44105.3 2
0
9 Inverter~
13 1447 266 0 2 22
0 42 43
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U13F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
6874 0 0
2
44105.3 1
0
14 Logic Display~
6 1450 232 0 1 2
10 43
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out43
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5305 0 0
2
44105.3 0
0
9 Inverter~
13 1401 266 0 2 22
0 44 45
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
34 0 0
2
44105.3 25
0
14 Logic Display~
6 1404 232 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out42
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
44105.3 24
0
9 Inverter~
13 1352 266 0 2 22
0 46 47
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
8402 0 0
2
44105.3 23
0
14 Logic Display~
6 1355 232 0 1 2
10 47
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out41
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3751 0 0
2
44105.3 22
0
9 Inverter~
13 1307 264 0 2 22
0 48 49
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
4292 0 0
2
44105.3 21
0
14 Logic Display~
6 1310 230 0 1 2
10 49
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out40
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6118 0 0
2
44105.3 20
0
9 Inverter~
13 1643 122 0 2 22
0 50 51
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
34 0 0
2
44105.3 19
0
14 Logic Display~
6 1646 88 0 1 2
10 51
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out39
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6357 0 0
2
44105.3 18
0
9 Inverter~
13 1596 114 0 2 22
0 63 52
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
319 0 0
2
44105.3 17
0
14 Logic Display~
6 1599 80 0 1 2
10 52
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out38
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3976 0 0
2
44105.3 16
0
9 Inverter~
13 1553 117 0 2 22
0 53 54
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U14F
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
7634 0 0
2
44105.3 15
0
14 Logic Display~
6 1556 83 0 1 2
10 54
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out37
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
523 0 0
2
44105.3 14
0
9 Inverter~
13 1502 119 0 2 22
0 55 56
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
6748 0 0
2
44105.3 13
0
14 Logic Display~
6 1505 85 0 1 2
10 56
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out36
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6901 0 0
2
44105.3 12
0
9 Inverter~
13 1448 118 0 2 22
0 57 58
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
842 0 0
2
44105.3 11
0
14 Logic Display~
6 1451 84 0 1 2
10 58
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Ou35
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3277 0 0
2
44105.3 10
0
9 Inverter~
13 1402 117 0 2 22
0 64 59
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
4212 0 0
2
44105.3 9
0
14 Logic Display~
6 1405 83 0 1 2
10 59
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out34
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4720 0 0
2
44105.3 8
0
9 Inverter~
13 1353 119 0 2 22
0 65 60
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
5551 0 0
2
44105.3 7
0
14 Logic Display~
6 1356 85 0 1 2
10 60
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out33
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6986 0 0
2
44105.3 6
0
14 Logic Display~
6 1310 85 0 1 2
10 61
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out32
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8745 0 0
2
44105.3 5
0
9 Inverter~
13 1307 119 0 2 22
0 62 61
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U15E
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 11 0
1 U
9592 0 0
2
44105.3 4
0
7 74LS138
19 1238 182 0 14 29
0 136 137 138 139 140 141 50 63 53
55 57 64 65 62
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U16
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 0 0 0 0
1 U
8748 0 0
2
44105.3 3
0
7 74LS138
19 1240 596 0 14 29
0 142 143 144 145 146 147 2 4 6
8 10 12 14 16
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U17
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 0 0 0 0
1 U
7168 0 0
2
44105.3 2
0
7 74LS138
19 1236 458 0 14 29
0 148 149 150 151 152 153 18 20 22
24 26 28 30 32
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U18
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 0 0 0 0
1 U
631 0 0
2
44105.3 1
0
7 74LS138
19 1237 328 0 14 29
0 154 155 156 157 158 159 34 36 38
40 42 44 46 48
0
0 0 5104 0
6 74F138
-21 -61 21 -53
3 U19
-10 -71 11 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 0 0 0 0
1 U
9466 0 0
2
44105.3 0
0
9 Inverter~
13 740 549 0 2 22
0 69 70
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
3266 0 0
2
44105.3 1
0
14 Logic Display~
6 743 515 0 1 2
10 70
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out31
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7693 0 0
2
44105.3 0
0
9 Inverter~
13 693 548 0 2 22
0 71 72
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
3723 0 0
2
44105.3 1
0
14 Logic Display~
6 696 514 0 1 2
10 72
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out30
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3440 0 0
2
44105.3 0
0
9 Inverter~
13 648 549 0 2 22
0 73 74
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U10A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
6263 0 0
2
44105.3 1
0
14 Logic Display~
6 651 515 0 1 2
10 74
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out29
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4900 0 0
2
44105.3 0
0
9 Inverter~
13 598 551 0 2 22
0 75 76
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 5 0
1 U
8783 0 0
2
44105.3 1
0
14 Logic Display~
6 601 517 0 1 2
10 76
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out28
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3221 0 0
2
44105.3 0
0
9 Inverter~
13 544 548 0 2 22
0 77 78
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 5 0
1 U
3215 0 0
2
44105.3 1
0
14 Logic Display~
6 547 514 0 1 2
10 78
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out27
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7903 0 0
2
44105.3 0
0
9 Inverter~
13 498 549 0 2 22
0 79 80
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
7121 0 0
2
44105.3 1
0
14 Logic Display~
6 501 515 0 1 2
10 80
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out26
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4484 0 0
2
44105.3 0
0
9 Inverter~
13 449 548 0 2 22
0 81 82
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
5996 0 0
2
44105.3 1
0
14 Logic Display~
6 452 514 0 1 2
10 82
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out25
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7804 0 0
2
44105.3 0
0
9 Inverter~
13 406 546 0 2 22
0 83 84
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
5523 0 0
2
44105.3 1
0
14 Logic Display~
6 409 512 0 1 2
10 84
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out24
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3330 0 0
2
44105.3 0
0
9 Inverter~
13 740 412 0 2 22
0 85 86
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U9A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3465 0 0
2
44105.3 1
0
14 Logic Display~
6 743 378 0 1 2
10 86
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out23
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8396 0 0
2
44105.3 0
0
9 Inverter~
13 693 411 0 2 22
0 87 88
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
3685 0 0
2
44105.3 1
0
14 Logic Display~
6 696 377 0 1 2
10 88
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out22
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7849 0 0
2
44105.3 0
0
9 Inverter~
13 650 410 0 2 22
0 89 90
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
6343 0 0
2
44105.3 1
0
14 Logic Display~
6 653 376 0 1 2
10 90
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out21
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7376 0 0
2
44105.3 0
0
9 Inverter~
13 599 412 0 2 22
0 91 92
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
9156 0 0
2
44105.3 1
0
14 Logic Display~
6 602 378 0 1 2
10 92
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out20
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5776 0 0
2
44105.3 0
0
9 Inverter~
13 545 413 0 2 22
0 93 94
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
7207 0 0
2
44105.3 1
0
14 Logic Display~
6 548 379 0 1 2
10 94
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out19
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4459 0 0
2
44105.3 0
0
9 Inverter~
13 499 412 0 2 22
0 95 96
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
3760 0 0
2
44105.3 1
0
14 Logic Display~
6 502 378 0 1 2
10 96
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out18
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
754 0 0
2
44105.3 0
0
9 Inverter~
13 450 412 0 2 22
0 97 98
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U8A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
9767 0 0
2
44105.3 1
0
14 Logic Display~
6 453 378 0 1 2
10 98
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out17
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7978 0 0
2
44105.3 0
0
9 Inverter~
13 407 413 0 2 22
0 99 100
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
3142 0 0
2
44105.3 1
0
14 Logic Display~
6 410 379 0 1 2
10 100
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out16
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3284 0 0
2
44105.3 0
0
9 Inverter~
13 736 276 0 2 22
0 101 102
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
659 0 0
2
44105.3 1
0
14 Logic Display~
6 739 242 0 1 2
10 102
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out15
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3800 0 0
2
44105.3 0
0
9 Inverter~
13 689 274 0 2 22
0 103 104
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
6792 0 0
2
44105.3 1
0
14 Logic Display~
6 692 240 0 1 2
10 104
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out14
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3701 0 0
2
44105.3 0
0
9 Inverter~
13 646 274 0 2 22
0 105 106
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
6316 0 0
2
44105.3 1
0
14 Logic Display~
6 649 240 0 1 2
10 106
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out13
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8734 0 0
2
44105.3 0
0
9 Inverter~
13 595 275 0 2 22
0 107 108
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
7988 0 0
2
44105.3 1
0
14 Logic Display~
6 598 241 0 1 2
10 108
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out12
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3217 0 0
2
44105.3 0
0
9 Inverter~
13 541 273 0 2 22
0 109 110
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3965 0 0
2
44105.3 1
0
14 Logic Display~
6 544 239 0 1 2
10 110
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out11
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8239 0 0
2
44105.3 0
0
9 Inverter~
13 495 273 0 2 22
0 111 112
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
828 0 0
2
44105.3 1
0
14 Logic Display~
6 498 239 0 1 2
10 112
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out10
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6187 0 0
2
44105.3 0
0
9 Inverter~
13 446 273 0 2 22
0 113 114
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
7107 0 0
2
44105.3 1
0
14 Logic Display~
6 449 239 0 1 2
10 114
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out9
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6433 0 0
2
44105.3 0
0
9 Inverter~
13 401 271 0 2 22
0 115 116
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
8559 0 0
2
44105.3 1
0
14 Logic Display~
6 404 237 0 1 2
10 116
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out8
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3674 0 0
2
44105.3 0
0
9 Inverter~
13 737 129 0 2 22
0 117 118
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
5697 0 0
2
44105.3 1
0
14 Logic Display~
6 740 95 0 1 2
10 118
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out7
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3805 0 0
2
44105.3 0
0
9 Inverter~
13 690 121 0 2 22
0 133 119
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
5219 0 0
2
44105.3 1
0
14 Logic Display~
6 693 87 0 1 2
10 119
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out6
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3795 0 0
2
44105.3 0
0
9 Inverter~
13 647 124 0 2 22
0 120 121
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3637 0 0
2
44105.3 1
0
14 Logic Display~
6 650 90 0 1 2
10 121
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out5
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3226 0 0
2
44105.3 0
0
9 Inverter~
13 596 126 0 2 22
0 122 123
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
6966 0 0
2
44105.3 1
0
14 Logic Display~
6 599 92 0 1 2
10 123
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out4
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9796 0 0
2
44105.3 0
0
9 Inverter~
13 542 125 0 2 22
0 124 125
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5952 0 0
2
44105.3 1
0
14 Logic Display~
6 545 91 0 1 2
10 125
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out3
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3649 0 0
2
44105.3 0
0
9 Inverter~
13 496 124 0 2 22
0 134 126
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3716 0 0
2
44105.3 1
0
14 Logic Display~
6 499 90 0 1 2
10 126
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out2
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4797 0 0
2
44105.3 0
0
9 Inverter~
13 447 126 0 2 22
0 135 127
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4681 0 0
2
44105.3 1
0
14 Logic Display~
6 450 92 0 1 2
10 127
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Out1
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9730 0 0
2
44105.3 0
0
14 Logic Display~
6 404 92 0 1 2
10 128
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 Out00
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9874 0 0
2
44105.3 0
0
9 Inverter~
13 401 126 0 2 22
0 129 128
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
364 0 0
2
44105.3 0
0
9 Inverter~
13 69 345 0 2 22
0 66 130
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3656 0 0
2
44105.3 0
0
7 74LS138
19 332 189 0 14 29
0 132 131 68 130 66 67 117 133 120
122 124 134 135 129
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
3131 0 0
2
44105.3 8
0
7 74LS138
19 334 603 0 14 29
0 132 131 68 67 130 130 69 71 73
75 77 79 81 83
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U4
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
6772 0 0
2
44105.3 0
0
7 74LS138
19 330 465 0 14 29
0 132 131 68 67 66 66 85 87 89
91 93 95 97 99
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U3
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
9557 0 0
2
44105.3 0
0
7 74LS138
19 331 335 0 14 29
0 132 131 68 66 67 67 101 103 105
107 109 111 113 115
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U2
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
5789 0 0
2
44105.3 8
0
209
1 0 2 0 0 4112 0 6 0 0 70 2
1649 560
1648 560
1 2 3 0 0 4240 0 7 6 0 0 2
1649 526
1649 524
1 0 4 0 0 4112 0 8 0 0 71 2
1602 559
1601 559
1 2 5 0 0 4240 0 9 8 0 0 2
1602 525
1602 523
1 0 6 0 0 4112 0 10 0 0 62 2
1557 560
1558 560
1 2 7 0 0 4240 0 11 10 0 0 2
1557 526
1557 524
1 0 8 0 0 16 0 12 0 0 72 2
1507 562
1507 562
1 2 9 0 0 4240 0 13 12 0 0 2
1507 528
1507 526
1 0 10 0 0 16 0 14 0 0 73 2
1453 559
1453 559
1 2 11 0 0 4240 0 15 14 0 0 2
1453 525
1453 523
1 0 12 0 0 16 0 16 0 0 74 2
1407 560
1407 560
1 2 13 0 0 4240 0 17 16 0 0 2
1407 526
1407 524
1 0 14 0 0 16 0 18 0 0 75 2
1358 559
1358 559
1 2 15 0 0 4240 0 19 18 0 0 2
1358 525
1358 523
1 0 16 0 0 16 0 20 0 0 76 2
1315 557
1315 557
1 2 17 0 0 4240 0 21 20 0 0 2
1315 523
1315 521
1 0 18 0 0 16 0 22 0 0 77 2
1649 423
1649 423
1 2 19 0 0 4240 0 23 22 0 0 2
1649 389
1649 387
1 0 20 0 0 16 0 24 0 0 78 2
1602 422
1602 422
1 2 21 0 0 4240 0 25 24 0 0 2
1602 388
1602 386
1 0 22 0 0 16 0 26 0 0 79 2
1559 421
1559 421
1 2 23 0 0 4240 0 27 26 0 0 2
1559 387
1559 385
1 0 24 0 0 16 0 28 0 0 80 2
1508 423
1508 423
1 2 25 0 0 4240 0 29 28 0 0 2
1508 389
1508 387
1 0 26 0 0 16 0 30 0 0 81 2
1454 424
1454 424
1 2 27 0 0 4240 0 31 30 0 0 2
1454 390
1454 388
1 0 28 0 0 16 0 32 0 0 82 2
1408 423
1408 423
1 2 29 0 0 4240 0 33 32 0 0 2
1408 389
1408 387
1 0 30 0 0 16 0 34 0 0 83 2
1359 423
1359 423
1 2 31 0 0 4240 0 35 34 0 0 2
1359 389
1359 387
1 0 32 0 0 16 0 36 0 0 84 2
1316 424
1316 424
1 2 33 0 0 4240 0 37 36 0 0 2
1316 390
1316 388
1 0 34 0 0 16 0 38 0 0 85 2
1645 287
1645 287
1 2 35 0 0 4240 0 39 38 0 0 2
1645 253
1645 251
1 0 36 0 0 16 0 40 0 0 86 2
1598 285
1598 285
1 2 37 0 0 4240 0 41 40 0 0 2
1598 251
1598 249
1 0 38 0 0 16 0 42 0 0 87 2
1555 285
1555 285
1 2 39 0 0 4240 0 43 42 0 0 2
1555 251
1555 249
1 0 40 0 0 16 0 44 0 0 88 2
1504 286
1504 286
1 2 41 0 0 4240 0 45 44 0 0 2
1504 252
1504 250
1 0 42 0 0 16 0 46 0 0 89 2
1450 284
1450 284
1 2 43 0 0 4240 0 47 46 0 0 2
1450 250
1450 248
1 0 44 0 0 16 0 48 0 0 90 2
1404 284
1404 284
1 2 45 0 0 4240 0 49 48 0 0 2
1404 250
1404 248
1 0 46 0 0 16 0 50 0 0 91 2
1355 284
1355 284
1 2 47 0 0 4240 0 51 50 0 0 2
1355 250
1355 248
1 0 48 0 0 16 0 52 0 0 92 2
1310 282
1310 282
1 2 49 0 0 4240 0 53 52 0 0 2
1310 248
1310 246
1 0 50 0 0 16 0 54 0 0 63 2
1646 140
1646 140
1 2 51 0 0 4240 0 55 54 0 0 2
1646 106
1646 104
1 2 52 0 0 4240 0 57 56 0 0 2
1599 98
1599 96
1 0 53 0 0 16 0 58 0 0 65 2
1556 135
1556 135
1 2 54 0 0 4240 0 59 58 0 0 2
1556 101
1556 99
1 0 55 0 0 16 0 60 0 0 66 2
1505 137
1505 137
1 2 56 0 0 4240 0 61 60 0 0 2
1505 103
1505 101
1 0 57 0 0 16 0 62 0 0 67 2
1451 136
1451 136
1 2 58 0 0 4240 0 63 62 0 0 2
1451 102
1451 100
1 2 59 0 0 4240 0 65 64 0 0 2
1405 101
1405 99
1 2 60 0 0 4240 0 67 66 0 0 2
1356 103
1356 101
1 2 61 0 0 4240 0 68 69 0 0 2
1310 103
1310 101
14 1 62 0 0 8336 0 70 69 0 0 3
1276 218
1310 218
1310 137
0 9 6 0 0 8336 0 0 71 0 0 3
1558 547
1558 587
1278 587
7 0 50 0 0 4240 0 70 0 0 0 3
1276 155
1646 155
1646 136
1 8 63 0 0 8336 0 56 70 0 0 3
1599 132
1599 164
1276 164
9 0 53 0 0 4240 0 70 0 0 0 3
1276 173
1556 173
1556 131
10 0 55 0 0 4240 0 70 0 0 0 3
1276 182
1505 182
1505 133
11 0 57 0 0 4240 0 70 0 0 0 3
1276 191
1451 191
1451 133
12 1 64 0 0 4240 0 70 64 0 0 3
1276 200
1405 200
1405 135
13 1 65 0 0 4240 0 70 66 0 0 3
1276 209
1356 209
1356 137
7 0 2 0 0 4240 0 71 0 0 0 3
1278 569
1648 569
1648 550
0 8 4 0 0 8336 0 0 71 0 0 3
1601 545
1601 578
1278 578
10 0 8 0 0 4240 0 71 0 0 0 3
1278 596
1507 596
1507 547
11 0 10 0 0 4240 0 71 0 0 0 3
1278 605
1453 605
1453 547
12 0 12 0 0 4240 0 71 0 0 0 3
1278 614
1407 614
1407 547
13 0 14 0 0 4240 0 71 0 0 0 3
1278 623
1358 623
1358 549
0 14 16 0 0 4240 0 0 71 0 0 3
1315 548
1315 632
1278 632
7 0 18 0 0 4240 0 72 0 0 0 3
1274 431
1649 431
1649 418
0 8 20 0 0 8336 0 0 72 0 0 3
1602 413
1602 440
1274 440
9 0 22 0 0 4240 0 72 0 0 0 3
1274 449
1559 449
1559 413
10 0 24 0 0 4240 0 72 0 0 0 3
1274 458
1508 458
1508 415
11 0 26 0 0 4240 0 72 0 0 0 3
1274 467
1454 467
1454 415
12 0 28 0 0 4240 0 72 0 0 0 3
1274 476
1408 476
1408 415
13 0 30 0 0 4240 0 72 0 0 0 3
1274 485
1359 485
1359 417
0 14 32 0 0 4240 0 0 72 0 0 3
1316 416
1316 494
1274 494
7 0 34 0 0 4240 0 73 0 0 0 3
1275 301
1645 301
1645 282
0 8 36 0 0 8336 0 0 73 0 0 3
1598 277
1598 310
1275 310
9 0 38 0 0 4240 0 73 0 0 0 3
1275 319
1555 319
1555 277
10 0 40 0 0 4240 0 73 0 0 0 3
1275 328
1504 328
1504 279
11 0 42 0 0 4240 0 73 0 0 0 3
1275 337
1450 337
1450 279
12 0 44 0 0 4240 0 73 0 0 0 3
1275 346
1404 346
1404 279
13 0 46 0 0 4240 0 73 0 0 0 3
1275 355
1355 355
1355 281
0 14 48 0 0 4240 0 0 73 0 0 3
1310 279
1310 364
1275 364
0 6 66 0 0 8192 0 0 141 94 0 3
140 492
140 501
292 501
0 5 66 0 0 8192 0 0 141 167 0 3
137 367
137 492
292 492
0 6 67 0 0 8192 0 0 142 163 0 3
153 372
153 371
293 371
0 5 67 0 0 0 0 0 142 163 0 3
153 364
153 362
293 362
0 3 68 0 0 8192 0 0 141 168 0 3
225 455
225 456
298 456
1 0 69 0 0 4096 0 74 0 0 187 2
743 567
742 567
1 2 70 0 0 4224 0 75 74 0 0 2
743 533
743 531
1 0 71 0 0 4096 0 76 0 0 188 2
696 566
695 566
1 2 72 0 0 4224 0 77 76 0 0 2
696 532
696 530
1 0 73 0 0 4096 0 78 0 0 179 2
651 567
652 567
1 2 74 0 0 4224 0 79 78 0 0 2
651 533
651 531
1 0 75 0 0 0 0 80 0 0 189 2
601 569
601 569
1 2 76 0 0 4224 0 81 80 0 0 2
601 535
601 533
1 0 77 0 0 0 0 82 0 0 190 2
547 566
547 566
1 2 78 0 0 4224 0 83 82 0 0 2
547 532
547 530
1 0 79 0 0 0 0 84 0 0 191 2
501 567
501 567
1 2 80 0 0 4224 0 85 84 0 0 2
501 533
501 531
1 0 81 0 0 0 0 86 0 0 192 2
452 566
452 566
1 2 82 0 0 4224 0 87 86 0 0 2
452 532
452 530
1 0 83 0 0 0 0 88 0 0 193 2
409 564
409 564
1 2 84 0 0 4224 0 89 88 0 0 2
409 530
409 528
1 0 85 0 0 0 0 90 0 0 194 2
743 430
743 430
1 2 86 0 0 4224 0 91 90 0 0 2
743 396
743 394
1 0 87 0 0 0 0 92 0 0 195 2
696 429
696 429
1 2 88 0 0 4224 0 93 92 0 0 2
696 395
696 393
1 0 89 0 0 0 0 94 0 0 196 2
653 428
653 428
1 2 90 0 0 4224 0 95 94 0 0 2
653 394
653 392
1 0 91 0 0 0 0 96 0 0 197 2
602 430
602 430
1 2 92 0 0 4224 0 97 96 0 0 2
602 396
602 394
1 0 93 0 0 0 0 98 0 0 198 2
548 431
548 431
1 2 94 0 0 4224 0 99 98 0 0 2
548 397
548 395
1 0 95 0 0 0 0 100 0 0 199 2
502 430
502 430
1 2 96 0 0 4224 0 101 100 0 0 2
502 396
502 394
1 0 97 0 0 0 0 102 0 0 200 2
453 430
453 430
1 2 98 0 0 4224 0 103 102 0 0 2
453 396
453 394
1 0 99 0 0 0 0 104 0 0 201 2
410 431
410 431
1 2 100 0 0 4224 0 105 104 0 0 2
410 397
410 395
1 0 101 0 0 0 0 106 0 0 202 2
739 294
739 294
1 2 102 0 0 4224 0 107 106 0 0 2
739 260
739 258
1 0 103 0 0 0 0 108 0 0 203 2
692 292
692 292
1 2 104 0 0 4224 0 109 108 0 0 2
692 258
692 256
1 0 105 0 0 0 0 110 0 0 204 2
649 292
649 292
1 2 106 0 0 4224 0 111 110 0 0 2
649 258
649 256
1 0 107 0 0 0 0 112 0 0 205 2
598 293
598 293
1 2 108 0 0 4224 0 113 112 0 0 2
598 259
598 257
1 0 109 0 0 0 0 114 0 0 206 2
544 291
544 291
1 2 110 0 0 4224 0 115 114 0 0 2
544 257
544 255
1 0 111 0 0 0 0 116 0 0 207 2
498 291
498 291
1 2 112 0 0 4224 0 117 116 0 0 2
498 257
498 255
1 0 113 0 0 0 0 118 0 0 208 2
449 291
449 291
1 2 114 0 0 4224 0 119 118 0 0 2
449 257
449 255
1 0 115 0 0 0 0 120 0 0 209 2
404 289
404 289
1 2 116 0 0 4224 0 121 120 0 0 2
404 255
404 253
1 0 117 0 0 0 0 122 0 0 180 2
740 147
740 147
1 2 118 0 0 4224 0 123 122 0 0 2
740 113
740 111
1 2 119 0 0 4224 0 125 124 0 0 2
693 105
693 103
1 0 120 0 0 0 0 126 0 0 182 2
650 142
650 142
1 2 121 0 0 4224 0 127 126 0 0 2
650 108
650 106
1 0 122 0 0 0 0 128 0 0 183 2
599 144
599 144
1 2 123 0 0 4224 0 129 128 0 0 2
599 110
599 108
1 0 124 0 0 0 0 130 0 0 184 2
545 143
545 143
1 2 125 0 0 4224 0 131 130 0 0 2
545 109
545 107
1 2 126 0 0 4224 0 133 132 0 0 2
499 108
499 106
1 2 127 0 0 4224 0 135 134 0 0 2
450 110
450 108
1 2 128 0 0 4224 0 136 137 0 0 2
404 110
404 108
14 1 129 0 0 8320 0 139 137 0 0 3
370 225
404 225
404 144
0 4 67 0 0 8192 0 0 140 162 0 3
153 483
153 621
302 621
0 6 130 0 0 8192 0 0 140 161 0 3
123 630
123 639
296 639
0 5 130 0 0 4224 0 0 140 165 0 3
123 345
123 630
296 630
0 4 67 0 0 0 0 0 141 163 0 3
153 411
153 483
298 483
1 6 67 0 0 8320 0 1 139 0 0 4
45 411
153 411
153 225
294 225
0 5 66 0 0 8192 0 0 139 167 0 3
138 354
138 216
294 216
2 4 130 0 0 0 0 138 139 0 0 4
90 345
124 345
124 207
300 207
0 1 66 0 0 0 0 0 138 167 0 2
54 367
54 345
1 4 66 0 0 12416 0 2 142 0 0 4
44 367
138 367
138 353
299 353
0 3 68 0 0 4224 0 0 140 169 0 3
225 326
225 594
302 594
0 3 68 0 0 0 0 0 142 176 0 3
225 180
225 326
299 326
0 2 131 0 0 4096 0 0 140 171 0 3
246 446
246 585
302 585
0 2 131 0 0 0 0 0 141 172 0 3
246 317
246 447
298 447
0 2 131 0 0 4096 0 0 142 177 0 3
246 171
246 317
299 317
0 1 132 0 0 4096 0 0 140 174 0 3
267 438
267 576
302 576
0 1 132 0 0 0 0 0 141 175 0 3
267 308
267 438
298 438
0 1 132 0 0 4096 0 0 142 178 0 3
267 162
267 308
299 308
1 3 68 0 0 0 0 5 139 0 0 4
75 263
95 263
95 180
300 180
1 2 131 0 0 12416 0 4 139 0 0 4
78 214
85 214
85 171
300 171
1 1 132 0 0 8320 0 3 139 0 0 3
79 163
79 162
300 162
0 9 73 0 0 8320 0 0 140 0 0 3
652 554
652 594
372 594
7 0 117 0 0 4224 0 139 0 0 0 3
370 162
740 162
740 143
1 8 133 0 0 8320 0 124 139 0 0 3
693 139
693 171
370 171
9 0 120 0 0 4224 0 139 0 0 0 3
370 180
650 180
650 138
10 0 122 0 0 4224 0 139 0 0 0 3
370 189
599 189
599 140
11 0 124 0 0 4224 0 139 0 0 0 3
370 198
545 198
545 140
12 1 134 0 0 4224 0 139 132 0 0 3
370 207
499 207
499 142
13 1 135 0 0 4224 0 139 134 0 0 3
370 216
450 216
450 144
7 0 69 0 0 4224 0 140 0 0 0 3
372 576
742 576
742 557
0 8 71 0 0 8320 0 0 140 0 0 3
695 552
695 585
372 585
10 0 75 0 0 4224 0 140 0 0 0 3
372 603
601 603
601 554
11 0 77 0 0 4224 0 140 0 0 0 3
372 612
547 612
547 554
12 0 79 0 0 4224 0 140 0 0 0 3
372 621
501 621
501 554
13 0 81 0 0 4224 0 140 0 0 0 3
372 630
452 630
452 556
0 14 83 0 0 4224 0 0 140 0 0 3
409 555
409 639
372 639
7 0 85 0 0 4224 0 141 0 0 0 3
368 438
743 438
743 425
0 8 87 0 0 8320 0 0 141 0 0 3
696 420
696 447
368 447
9 0 89 0 0 4224 0 141 0 0 0 3
368 456
653 456
653 420
10 0 91 0 0 4224 0 141 0 0 0 3
368 465
602 465
602 422
11 0 93 0 0 4224 0 141 0 0 0 3
368 474
548 474
548 422
12 0 95 0 0 4224 0 141 0 0 0 3
368 483
502 483
502 422
13 0 97 0 0 4224 0 141 0 0 0 3
368 492
453 492
453 424
0 14 99 0 0 4224 0 0 141 0 0 3
410 423
410 501
368 501
7 0 101 0 0 4224 0 142 0 0 0 3
369 308
739 308
739 289
0 8 103 0 0 8320 0 0 142 0 0 3
692 284
692 317
369 317
9 0 105 0 0 4224 0 142 0 0 0 3
369 326
649 326
649 284
10 0 107 0 0 4224 0 142 0 0 0 3
369 335
598 335
598 286
11 0 109 0 0 4224 0 142 0 0 0 3
369 344
544 344
544 286
12 0 111 0 0 4224 0 142 0 0 0 3
369 353
498 353
498 286
13 0 113 0 0 4224 0 142 0 0 0 3
369 362
449 362
449 288
0 14 115 0 0 4224 0 0 142 0 0 3
404 286
404 371
369 371
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
841 221 1022 245
851 229 1011 245
20 E=0 D=1, IC 2 active
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
840 191 949 215
850 199 938 215
11 Input 01011
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
841 248 934 272
851 256 923 272
9 Output 11
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
