CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 490 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
85
13 Logic Switch~
5 1062 498 0 1 11
0 14
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 S2
-2 -32 12 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3330 0 0
2
44087.4 0
0
13 Logic Switch~
5 1101 725 0 1 11
0 15
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 V0
-2 -29 12 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3465 0 0
2
44087.4 0
0
13 Logic Switch~
5 284 1403 0 1 11
0 26
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 B3
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8396 0 0
2
44087.4 10
0
13 Logic Switch~
5 266 1183 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-2 -18 12 -10
2 B2
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3685 0 0
2
44087.4 9
0
13 Logic Switch~
5 238 983 0 1 11
0 34
0
0 0 21360 0
2 0V
-2 -18 12 -10
2 B1
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7849 0 0
2
44087.4 8
0
13 Logic Switch~
5 232 756 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-2 -18 12 -10
2 B0
-3 -29 11 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6343 0 0
2
44087.4 7
0
13 Logic Switch~
5 552 875 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7376 0 0
2
44087.4 6
0
13 Logic Switch~
5 547 739 0 10 11
0 58 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9156 0 0
2
44087.4 5
0
13 Logic Switch~
5 556 957 0 10 11
0 53 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5776 0 0
2
44087.4 4
0
13 Logic Switch~
5 545 1165 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7207 0 0
2
44087.4 3
0
13 Logic Switch~
5 551 1380 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4459 0 0
2
44087.4 2
0
13 Logic Switch~
5 478 629 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S1
-10 -27 4 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3760 0 0
2
44087.4 35
0
13 Logic Switch~
5 430 694 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
754 0 0
2
44087.4 34
0
13 Logic Switch~
5 894 190 0 1 11
0 68
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9767 0 0
2
44087.4 33
0
13 Logic Switch~
5 588 81 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7978 0 0
2
44087.4 32
0
13 Logic Switch~
5 574 197 0 10 11
0 67 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3142 0 0
2
44087.4 31
0
13 Logic Switch~
5 572 501 0 1 11
0 65
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3284 0 0
2
44087.4 30
0
13 Logic Switch~
5 586 385 0 1 11
0 64
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
659 0 0
2
44087.4 29
0
13 Logic Switch~
5 884 375 0 1 11
0 59
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3800 0 0
2
44087.4 28
0
13 Logic Switch~
5 396 374 0 1 11
0 73
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6792 0 0
2
44087.4 27
0
13 Logic Switch~
5 98 384 0 10 11
0 78 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3701 0 0
2
44087.4 26
0
13 Logic Switch~
5 84 500 0 1 11
0 79
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6316 0 0
2
44087.4 25
0
13 Logic Switch~
5 86 196 0 10 11
0 81 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8734 0 0
2
44087.4 24
0
13 Logic Switch~
5 100 80 0 10 11
0 80 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7988 0 0
2
44087.4 23
0
13 Logic Switch~
5 406 189 0 1 11
0 82
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3217 0 0
2
44087.4 22
0
14 Logic Display~
6 1391 559 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3965 0 0
2
44087.5 0
0
14 Logic Display~
6 1348 548 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8239 0 0
2
44087.5 0
0
14 Logic Display~
6 1313 544 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
828 0 0
2
44087.5 0
0
14 Logic Display~
6 1275 526 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Y3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6187 0 0
2
44087.5 0
0
7 74LS157
122 1223 593 0 14 29
0 14 9 5 8 4 7 3 6 2
15 13 12 11 10
0
0 0 4848 0
6 74F157
-21 -60 21 -52
3 U21
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
7107 0 0
2
44087.4 1
0
8 2-In OR~
219 452 1421 0 3 22
0 23 24 22
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U17B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
6433 0 0
2
44087.4 51
0
9 2-In AND~
219 386 1360 0 3 22
0 19 26 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
8559 0 0
2
44087.4 50
0
9 2-In AND~
219 388 1457 0 3 22
0 25 18 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3674 0 0
2
44087.4 49
0
9 Inverter~
13 327 1437 0 2 22
0 26 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
5697 0 0
2
44087.4 48
0
8 2-In OR~
219 436 1205 0 3 22
0 27 28 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U17A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3805 0 0
2
44087.4 47
0
9 2-In AND~
219 368 1140 0 3 22
0 19 30 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
5219 0 0
2
44087.4 46
0
9 2-In AND~
219 370 1237 0 3 22
0 29 18 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
3795 0 0
2
44087.4 45
0
9 Inverter~
13 309 1217 0 2 22
0 30 29
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
3637 0 0
2
44087.4 44
0
8 2-In OR~
219 414 997 0 3 22
0 31 32 52
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
3226 0 0
2
44087.4 43
0
9 2-In AND~
219 340 940 0 3 22
0 19 34 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6966 0 0
2
44087.4 42
0
9 2-In AND~
219 342 1037 0 3 22
0 33 18 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
9796 0 0
2
44087.4 41
0
9 Inverter~
13 281 1017 0 2 22
0 34 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
5952 0 0
2
44087.4 40
0
8 2-In OR~
219 407 779 0 3 22
0 35 36 57
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3649 0 0
2
44087.4 39
0
9 2-In AND~
219 334 713 0 3 22
0 19 38 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3716 0 0
2
44087.4 38
0
9 2-In AND~
219 336 810 0 3 22
0 37 18 36
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4797 0 0
2
44087.4 37
0
9 Inverter~
13 275 790 0 2 22
0 38 37
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
4681 0 0
2
44087.4 36
0
9 2-In XOR~
219 779 765 0 3 22
0 54 39 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9730 0 0
2
44087.4 34
0
9 2-In AND~
219 729 863 0 3 22
0 54 39 55
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9874 0 0
2
44087.4 33
0
8 2-In OR~
219 807 857 0 3 22
0 56 55 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
364 0 0
2
44087.4 32
0
9 2-In AND~
219 625 817 0 3 22
0 58 57 56
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3656 0 0
2
44087.4 31
0
9 2-In XOR~
219 656 756 0 3 22
0 58 57 54
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3131 0 0
2
44087.4 30
0
9 2-In XOR~
219 665 974 0 3 22
0 53 52 49
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
6772 0 0
2
44087.4 29
0
9 2-In AND~
219 634 1035 0 3 22
0 53 52 51
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9557 0 0
2
44087.4 28
0
8 2-In OR~
219 815 1072 0 3 22
0 51 50 16
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
5789 0 0
2
44087.4 27
0
9 2-In AND~
219 738 1081 0 3 22
0 49 20 50
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7328 0 0
2
44087.4 26
0
9 2-In XOR~
219 788 983 0 3 22
0 49 20 4
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4799 0 0
2
44087.4 25
0
9 2-In XOR~
219 654 1182 0 3 22
0 48 21 45
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9196 0 0
2
44087.4 23
0
9 2-In AND~
219 623 1243 0 3 22
0 48 21 47
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3857 0 0
2
44087.4 22
0
8 2-In OR~
219 805 1281 0 3 22
0 47 46 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7125 0 0
2
44087.4 21
0
9 2-In AND~
219 727 1290 0 3 22
0 45 16 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3641 0 0
2
44087.4 20
0
9 2-In XOR~
219 777 1191 0 3 22
0 45 16 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9821 0 0
2
44087.4 19
0
9 2-In XOR~
219 660 1397 0 3 22
0 44 22 41
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
3187 0 0
2
44087.4 17
0
9 2-In AND~
219 629 1458 0 3 22
0 44 22 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
762 0 0
2
44087.4 16
0
8 2-In OR~
219 810 1495 0 3 22
0 43 42 40
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
39 0 0
2
44087.4 15
0
9 2-In AND~
219 733 1504 0 3 22
0 41 17 42
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
9450 0 0
2
44087.4 14
0
9 2-In XOR~
219 783 1406 0 3 22
0 41 17 2
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3236 0 0
2
44087.4 13
0
14 Logic Display~
6 888 1477 0 1 2
10 40
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3321 0 0
2
44087.4 11
0
7 74LS153
119 852 274 0 14 29
0 72 71 70 69 18 19 63 60 62
61 68 59 7 6
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
8879 0 0
2
44087.4 21
0
9 2-In AND~
219 687 265 0 3 22
0 66 67 69
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
5433 0 0
2
44087.4 20
0
8 2-In OR~
219 683 188 0 3 22
0 66 67 70
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U17C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
3679 0 0
2
44087.4 19
0
9 2-In XOR~
219 688 134 0 3 22
0 66 67 71
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
9342 0 0
2
44087.4 18
0
9 Inverter~
13 686 81 0 2 22
0 66 72
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
3623 0 0
2
44087.4 17
0
9 Inverter~
13 684 385 0 2 22
0 64 63
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
3722 0 0
2
44087.4 15
0
9 2-In XOR~
219 688 439 0 3 22
0 64 65 60
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U10A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
8993 0 0
2
44087.4 14
0
8 2-In OR~
219 681 492 0 3 22
0 64 65 62
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U17D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
3723 0 0
2
44087.4 13
0
9 2-In AND~
219 690 543 0 3 22
0 64 65 61
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
6244 0 0
2
44087.4 12
0
9 2-In AND~
219 202 542 0 3 22
0 78 79 75
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
6421 0 0
2
44087.4 9
0
8 2-In OR~
219 193 491 0 3 22
0 78 79 76
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
7743 0 0
2
44087.4 8
0
9 2-In XOR~
219 200 438 0 3 22
0 78 79 74
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U10B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
9840 0 0
2
44087.4 7
0
9 Inverter~
13 196 384 0 2 22
0 78 77
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U15F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
6910 0 0
2
44087.4 6
0
9 Inverter~
13 198 80 0 2 22
0 80 86
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U13A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 17 0
1 U
449 0 0
2
44087.4 4
0
9 2-In XOR~
219 200 133 0 3 22
0 80 81 85
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U10C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
8761 0 0
2
44087.4 3
0
8 2-In OR~
219 195 187 0 3 22
0 80 81 84
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
6748 0 0
2
44087.4 2
0
9 2-In AND~
219 199 264 0 3 22
0 80 81 83
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U19A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
7393 0 0
2
44087.4 1
0
7 74LS153
119 365 268 0 14 29
0 86 85 84 83 18 19 77 74 76
75 82 73 9 8
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
3 U20
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 0 1 0 0 0
1 U
7699 0 0
2
44087.4 0
0
138
3 9 2 0 0 8320 0 66 30 0 0 4
816 1406
1125 1406
1125 629
1191 629
7 3 3 0 0 8320 0 30 61 0 0 4
1191 611
1068 611
1068 1191
810 1191
3 5 4 0 0 8320 0 56 30 0 0 4
821 983
1037 983
1037 593
1191 593
3 3 5 0 0 4224 0 30 47 0 0 4
1191 575
977 575
977 765
812 765
14 8 6 0 0 8320 0 68 30 0 0 4
884 301
1006 301
1006 620
1191 620
6 13 7 0 0 8320 0 30 68 0 0 4
1191 602
1123 602
1123 256
884 256
14 4 8 0 0 4224 0 85 30 0 0 4
397 295
1183 295
1183 584
1191 584
2 13 9 0 0 4224 0 30 85 0 0 4
1191 566
459 566
459 250
397 250
14 1 10 0 0 8320 0 30 29 0 0 3
1255 629
1275 629
1275 544
13 1 11 0 0 4224 0 30 28 0 0 3
1255 611
1313 611
1313 562
12 1 12 0 0 4240 0 30 27 0 0 4
1255 593
1334 593
1334 566
1348 566
11 1 13 0 0 12416 0 30 26 0 0 4
1255 575
1270 575
1270 577
1391 577
1 1 14 0 0 12416 0 1 30 0 0 4
1074 498
1097 498
1097 557
1191 557
1 10 15 0 0 8320 0 2 30 0 0 4
1113 725
1143 725
1143 638
1185 638
0 2 16 0 0 4096 0 0 61 16 0 3
673 1298
673 1200
761 1200
3 2 16 0 0 8320 0 54 60 0 0 7
848 1072
848 1140
567 1140
567 1298
673 1298
673 1299
703 1299
0 2 17 0 0 4096 0 0 65 53 0 2
667 1513
709 1513
0 2 18 0 0 8192 0 0 37 21 0 3
172 1248
172 1246
346 1246
0 2 18 0 0 4096 0 0 45 20 0 3
172 1048
172 819
312 819
0 2 18 0 0 0 0 0 41 21 0 3
172 1089
172 1046
318 1046
0 2 18 0 0 8320 0 0 33 87 0 6
489 570
62 570
62 1089
172 1089
172 1466
364 1466
1 0 19 0 0 4096 0 36 0 0 23 2
344 1131
126 1131
0 1 19 0 0 4224 0 0 32 25 0 3
126 969
126 1351
362 1351
1 0 19 0 0 0 0 40 0 0 25 2
316 931
126 931
1 0 19 0 0 0 0 44 0 0 89 6
310 704
126 704
126 971
91 971
91 598
442 598
0 2 20 0 0 4096 0 0 55 70 0 2
673 1090
714 1090
3 0 21 0 0 4224 0 35 0 0 67 2
469 1205
562 1205
3 0 22 0 0 8320 0 31 0 0 59 3
485 1421
485 1420
569 1420
3 1 23 0 0 4224 0 32 31 0 0 3
407 1360
407 1412
439 1412
3 2 24 0 0 8320 0 33 31 0 0 3
409 1457
409 1430
439 1430
2 1 25 0 0 8320 0 34 33 0 0 3
348 1437
348 1448
364 1448
1 2 26 0 0 4224 0 3 32 0 0 4
296 1403
337 1403
337 1369
362 1369
1 1 26 0 0 0 0 3 34 0 0 3
296 1403
296 1437
312 1437
3 1 27 0 0 4224 0 36 35 0 0 3
389 1140
389 1196
423 1196
3 2 28 0 0 8320 0 37 35 0 0 3
391 1237
391 1214
423 1214
2 1 29 0 0 8320 0 38 37 0 0 3
330 1217
330 1228
346 1228
1 2 30 0 0 4224 0 4 36 0 0 4
278 1183
319 1183
319 1149
344 1149
1 1 30 0 0 0 0 4 38 0 0 3
278 1183
278 1217
294 1217
3 1 31 0 0 4224 0 40 39 0 0 3
361 940
361 988
401 988
3 2 32 0 0 8320 0 41 39 0 0 3
363 1037
363 1006
401 1006
2 1 33 0 0 8320 0 42 41 0 0 3
302 1017
302 1028
318 1028
1 2 34 0 0 4224 0 5 40 0 0 4
250 983
291 983
291 949
316 949
1 1 34 0 0 0 0 5 42 0 0 3
250 983
250 1017
266 1017
3 1 35 0 0 4224 0 44 43 0 0 3
355 713
355 770
394 770
3 2 36 0 0 8320 0 45 43 0 0 3
357 810
357 788
394 788
2 1 37 0 0 8320 0 46 45 0 0 3
296 790
296 801
312 801
1 2 38 0 0 4224 0 6 44 0 0 4
244 756
285 756
285 722
310 722
1 1 38 0 0 0 0 6 46 0 0 3
244 756
244 790
260 790
0 2 39 0 0 4096 0 0 48 79 0 2
663 872
705 872
3 1 40 0 0 4224 0 0 67 51 0 2
865 1495
888 1495
3 0 40 0 0 0 0 64 0 0 50 2
843 1495
866 1495
0 1 41 0 0 4096 0 0 66 56 0 2
709 1397
767 1397
3 2 17 0 0 8320 0 59 66 0 0 7
838 1281
838 1339
564 1339
564 1513
668 1513
668 1415
767 1415
3 2 42 0 0 4224 0 65 64 0 0 2
754 1504
797 1504
3 1 43 0 0 4224 0 63 64 0 0 4
650 1458
767 1458
767 1486
797 1486
3 1 41 0 0 8320 0 62 65 0 0 3
693 1397
709 1397
709 1495
0 2 22 0 0 0 0 0 63 59 0 3
585 1420
585 1467
605 1467
0 1 44 0 0 4224 0 0 63 60 0 3
598 1380
598 1449
605 1449
0 2 22 0 0 0 0 0 62 0 0 4
564 1420
610 1420
610 1406
644 1406
1 1 44 0 0 0 0 11 62 0 0 4
563 1380
610 1380
610 1388
644 1388
0 1 45 0 0 4096 0 0 61 64 0 2
703 1182
761 1182
3 2 46 0 0 4224 0 60 59 0 0 2
748 1290
792 1290
3 1 47 0 0 4224 0 58 59 0 0 4
644 1243
761 1243
761 1272
792 1272
3 1 45 0 0 8320 0 57 60 0 0 3
687 1182
703 1182
703 1281
0 2 21 0 0 0 0 0 58 67 0 3
579 1205
579 1252
599 1252
0 1 48 0 0 4224 0 0 58 68 0 3
592 1165
592 1234
599 1234
0 2 21 0 0 0 0 0 57 0 0 4
558 1205
604 1205
604 1191
638 1191
1 1 48 0 0 0 0 10 57 0 0 4
557 1165
604 1165
604 1173
638 1173
0 1 49 0 0 4096 0 0 56 73 0 2
714 974
772 974
3 2 20 0 0 12416 0 49 56 0 0 8
840 857
868 857
868 913
577 913
577 1090
673 1090
673 992
772 992
3 2 50 0 0 4224 0 55 54 0 0 2
759 1081
802 1081
3 1 51 0 0 4224 0 53 54 0 0 4
655 1035
772 1035
772 1063
802 1063
3 1 49 0 0 8320 0 52 55 0 0 3
698 974
714 974
714 1072
0 2 52 0 0 4096 0 0 53 76 0 3
590 997
590 1044
610 1044
0 1 53 0 0 4224 0 0 53 77 0 3
603 957
603 1026
610 1026
3 2 52 0 0 4224 0 39 52 0 0 4
447 997
615 997
615 983
649 983
1 1 53 0 0 0 0 9 52 0 0 4
568 957
615 957
615 965
649 965
0 1 54 0 0 4096 0 0 47 82 0 2
705 756
763 756
1 2 39 0 0 8320 0 7 47 0 0 5
564 875
564 872
664 872
664 774
763 774
3 2 55 0 0 12416 0 48 49 0 0 4
750 863
765 863
765 866
794 866
3 1 56 0 0 4224 0 50 49 0 0 4
646 817
763 817
763 848
794 848
3 1 54 0 0 8320 0 51 48 0 0 3
689 756
705 756
705 854
0 2 57 0 0 4096 0 0 50 85 0 3
581 779
581 826
601 826
0 1 58 0 0 4224 0 0 50 86 0 3
594 739
594 808
601 808
3 2 57 0 0 4224 0 43 51 0 0 4
440 779
606 779
606 765
640 765
1 1 58 0 0 0 0 8 51 0 0 4
559 739
606 739
606 747
640 747
1 5 18 0 0 128 0 12 85 0 0 7
490 629
490 570
489 570
489 344
269 344
269 268
333 268
1 6 19 0 0 0 0 13 68 0 0 6
442 694
545 694
545 328
744 328
744 283
820 283
1 6 19 0 0 128 0 13 85 0 0 5
442 694
442 401
296 401
296 277
333 277
1 5 18 0 0 0 0 12 68 0 0 4
490 629
715 629
715 274
820 274
1 12 59 0 0 8320 0 19 68 0 0 4
896 375
910 375
910 319
890 319
8 3 60 0 0 8320 0 68 74 0 0 4
820 301
804 301
804 439
721 439
3 10 61 0 0 8320 0 76 68 0 0 3
711 543
820 543
820 319
3 9 62 0 0 8320 0 75 68 0 0 4
714 492
810 492
810 310
820 310
2 7 63 0 0 8320 0 73 68 0 0 4
705 385
797 385
797 292
820 292
0 1 64 0 0 4096 0 0 74 98 0 2
629 430
672 430
0 1 64 0 0 0 0 0 75 98 0 2
629 483
668 483
0 1 64 0 0 4224 0 0 76 99 0 3
629 385
629 534
666 534
1 1 64 0 0 0 0 18 73 0 0 2
598 385
669 385
1 2 65 0 0 8192 0 17 76 0 0 3
584 501
584 552
666 552
1 2 65 0 0 4096 0 17 75 0 0 2
584 501
668 501
1 2 65 0 0 8320 0 17 74 0 0 3
584 501
584 448
672 448
0 1 66 0 0 8192 0 0 71 105 0 3
631 126
631 125
672 125
0 1 66 0 0 0 0 0 70 105 0 2
631 179
670 179
0 1 66 0 0 4224 0 0 69 106 0 3
631 81
631 256
663 256
1 1 66 0 0 0 0 15 72 0 0 2
600 81
671 81
1 2 67 0 0 4096 0 16 69 0 0 3
586 197
586 274
663 274
1 2 67 0 0 4096 0 16 70 0 0 2
586 197
670 197
1 2 67 0 0 8320 0 16 71 0 0 3
586 197
586 143
672 143
1 11 68 0 0 4224 0 14 68 0 0 3
906 190
906 238
890 238
3 4 69 0 0 4224 0 69 68 0 0 2
708 265
820 265
3 3 70 0 0 12416 0 70 68 0 0 4
716 188
719 188
719 256
820 256
3 2 71 0 0 8320 0 71 68 0 0 4
721 134
728 134
728 247
820 247
2 1 72 0 0 8320 0 72 68 0 0 4
707 81
751 81
751 238
820 238
1 12 73 0 0 8320 0 20 85 0 0 4
408 374
422 374
422 313
403 313
8 3 74 0 0 8320 0 85 79 0 0 4
333 295
316 295
316 438
233 438
3 10 75 0 0 8320 0 77 85 0 0 3
223 542
333 542
333 313
3 9 76 0 0 8320 0 78 85 0 0 4
226 491
322 491
322 304
333 304
2 7 77 0 0 8320 0 80 85 0 0 4
217 384
309 384
309 286
333 286
0 1 78 0 0 4096 0 0 79 122 0 2
141 429
184 429
0 1 78 0 0 0 0 0 78 122 0 2
141 482
180 482
0 1 78 0 0 4224 0 0 77 123 0 3
141 384
141 533
178 533
1 1 78 0 0 0 0 21 80 0 0 2
110 384
181 384
1 2 79 0 0 8192 0 22 77 0 0 3
96 500
96 551
178 551
1 2 79 0 0 4096 0 22 78 0 0 2
96 500
180 500
1 2 79 0 0 8320 0 22 79 0 0 3
96 500
96 447
184 447
0 1 80 0 0 8192 0 0 82 129 0 3
143 125
143 124
184 124
0 1 80 0 0 0 0 0 83 129 0 2
143 178
182 178
0 1 80 0 0 4224 0 0 84 130 0 3
143 80
143 255
175 255
1 1 80 0 0 0 0 24 81 0 0 2
112 80
183 80
1 2 81 0 0 4096 0 23 84 0 0 3
98 196
98 273
175 273
1 2 81 0 0 4096 0 23 83 0 0 2
98 196
182 196
1 2 81 0 0 8320 0 23 82 0 0 3
98 196
98 142
184 142
1 11 82 0 0 4224 0 25 85 0 0 3
418 189
418 232
403 232
3 4 83 0 0 12416 0 84 85 0 0 4
220 264
235 264
235 259
333 259
3 3 84 0 0 12416 0 83 85 0 0 4
228 187
231 187
231 250
333 250
3 2 85 0 0 8320 0 82 85 0 0 4
233 133
240 133
240 241
333 241
2 1 86 0 0 8320 0 81 85 0 0 4
219 80
263 80
263 232
333 232
109
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
940 1411 971 1435
949 1420 961 1436
2 Y3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
928 1198 959 1222
937 1207 949 1223
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
939 991 970 1015
948 1000 960 1016
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
920 771 951 795
929 780 941 796
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
743 1500 770 1524
748 1505 764 1521
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
698 1516 725 1540
703 1521 719 1537
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
688 1478 715 1502
693 1483 709 1499
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
643 1436 664 1460
649 1441 657 1457
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
594 1468 613 1492
599 1473 607 1489
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
594 1421 621 1445
599 1427 615 1443
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
805 1405 834 1429
811 1411 827 1427
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
753 1418 780 1442
758 1423 774 1439
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
753 1368 782 1392
759 1373 775 1389
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
683 1375 706 1399
690 1381 698 1397
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
631 1355 660 1379
637 1361 653 1377
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
688 949 711 973
695 955 703 971
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
637 933 664 957
642 939 658 955
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
809 982 840 1006
816 987 832 1003
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
755 944 786 968
762 949 778 965
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
635 1408 656 1432
641 1413 649 1429
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
835 1473 862 1497
840 1479 856 1495
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
781 1509 810 1533
787 1515 803 1531
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
780 1462 807 1486
785 1467 801 1483
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
832 1258 851 1282
837 1263 845 1279
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
778 1294 797 1318
783 1299 791 1315
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
774 1247 801 1271
779 1253 795 1269
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
843 1050 862 1074
848 1055 856 1071
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
787 1087 808 1111
793 1093 801 1109
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
785 1040 806 1064
791 1045 799 1061
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
749 1080 776 1104
754 1085 770 1101
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
699 1094 726 1118
704 1099 720 1115
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
695 1053 722 1077
700 1058 716 1074
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
648 1013 667 1037
653 1019 661 1035
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
597 1045 616 1069
602 1050 610 1066
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
597 998 624 1022
602 1003 618 1019
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
757 995 786 1019
763 1001 779 1017
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
640 985 659 1009
645 991 653 1007
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
897 1488 944 1512
904 1494 936 1510
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
628 1141 649 1165
634 1147 642 1163
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
590 1206 611 1230
596 1212 604 1228
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
629 1193 648 1217
634 1198 642 1214
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
588 1253 607 1277
593 1258 601 1274
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
680 1158 699 1182
685 1163 693 1179
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
637 1221 656 1245
642 1226 650 1242
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
751 1152 770 1176
756 1158 764 1174
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
687 1259 706 1283
692 1265 700 1281
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
692 1301 713 1325
698 1306 706 1322
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
741 1285 760 1309
746 1291 754 1307
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
751 1203 772 1227
757 1208 765 1224
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
802 1190 821 1214
807 1196 815 1212
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
804 764 823 788
809 770 817 786
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
753 777 774 801
759 782 767 798
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
743 859 762 883
748 865 756 881
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
694 875 715 899
700 880 708 896
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
689 833 708 857
694 839 702 855
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
753 726 772 750
758 732 766 748
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
639 795 658 819
644 800 652 816
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
834 832 853 856
839 837 847 853
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
682 732 701 756
687 737 695 753
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
780 868 799 892
785 873 793 889
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
590 827 609 851
595 832 603 848
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
631 767 650 791
636 772 644 788
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
779 821 800 845
785 827 793 843
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
592 780 613 804
598 786 606 802
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
630 715 651 739
636 721 644 737
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
712 411 747 433
721 418 737 434
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
705 466 740 488
714 473 730 489
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
700 518 735 540
709 525 725 541
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
647 554 682 576
656 561 672 577
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
646 496 681 518
655 503 671 519
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
651 441 686 463
660 448 676 464
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
641 510 676 532
650 517 666 533
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
642 457 677 479
651 464 667 480
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
647 404 682 426
656 411 672 427
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
708 110 733 132
716 117 724 133
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
701 165 726 187
709 172 717 188
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
698 246 723 268
706 253 714 269
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
695 359 720 381
703 366 711 382
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
651 357 678 379
660 365 668 381
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
648 269 675 291
657 277 665 293
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
650 196 677 218
659 204 667 220
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
648 137 675 159
657 145 665 161
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
645 234 678 256
653 241 669 257
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
644 156 677 178
652 163 668 179
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
645 99 678 121
653 106 669 122
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
214 520 237 542
221 528 229 544
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
218 465 241 487
225 473 233 489
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
224 413 247 435
231 421 239 437
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
699 57 722 79
706 65 714 81
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
653 53 678 75
661 60 669 76
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
166 551 191 573
174 558 182 574
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
167 496 192 518
175 504 183 520
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
166 442 191 464
174 449 182 465
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
165 511 190 533
173 519 181 535
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
171 453 196 475
179 461 187 477
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
167 404 192 426
175 412 183 428
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
207 357 232 379
215 365 223 381
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
226 111 251 133
234 118 242 134
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
217 165 242 187
225 172 233 188
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
217 268 242 290
225 275 233 291
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
162 358 187 380
170 365 178 381
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
213 55 236 77
220 63 228 79
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
174 137 197 159
181 145 189 161
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
168 199 191 221
175 207 183 223
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
164 276 187 298
171 284 179 300
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
164 225 191 247
173 233 181 249
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
165 149 192 171
174 157 182 173
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
169 94 196 116
178 102 186 118
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
166 51 193 73
175 59 183 75
1 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
