CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
109
13 Logic Switch~
5 75 217 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S1
-8 -26 6 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44059.4 0
0
13 Logic Switch~
5 84 90 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44059.4 0
0
13 Logic Switch~
5 311 257 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44059.4 8
0
13 Logic Switch~
5 306 121 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44059.4 7
0
13 Logic Switch~
5 835 179 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44059.4 8
0
13 Logic Switch~
5 836 138 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44059.4 7
0
13 Logic Switch~
5 866 49 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
44059.4 6
0
13 Logic Switch~
5 846 343 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-5 -27 9 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44059.4 5
0
13 Logic Switch~
5 842 296 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
44059.4 4
0
13 Logic Switch~
5 840 253 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
44059.4 3
0
13 Logic Switch~
5 860 215 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
44059.4 2
0
13 Logic Switch~
5 949 373 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 Cin1
-12 -26 16 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
44059.4 1
0
13 Logic Switch~
5 845 92 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
44059.4 0
0
13 Logic Switch~
5 29 142 0 1 11
0 7
0
0 0 21360 0
2 0V
-2 -18 12 -10
1 B
0 -29 7 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
44059.4 0
0
13 Logic Switch~
5 191 1353 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3835 0 0
2
44059.4 1
0
13 Logic Switch~
5 191 1403 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
44059.4 0
0
13 Logic Switch~
5 756 967 0 1 11
0 49
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.89948e-315 5.38788e-315
0
13 Logic Switch~
5 616 1348 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
4 Cin3
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9323 0 0
2
5.89948e-315 5.37752e-315
0
13 Logic Switch~
5 625 1090 0 1 11
0 40
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.89948e-315 5.36716e-315
0
13 Logic Switch~
5 623 1138 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -16 7 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3108 0 0
2
5.89948e-315 5.3568e-315
0
13 Logic Switch~
5 615 1199 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4299 0 0
2
5.89948e-315 5.34643e-315
0
13 Logic Switch~
5 618 1269 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-5 -30 9 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9672 0 0
2
5.89948e-315 5.32571e-315
0
13 Logic Switch~
5 777 924 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7876 0 0
2
5.89948e-315 5.30499e-315
0
13 Logic Switch~
5 747 1013 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
5.89948e-315 5.26354e-315
0
13 Logic Switch~
5 746 1054 0 1 11
0 51
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.89948e-315 0
0
13 Logic Switch~
5 761 591 0 1 11
0 69
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
5.89948e-315 5.38788e-315
0
13 Logic Switch~
5 762 550 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3820 0 0
2
5.89948e-315 5.37752e-315
0
13 Logic Switch~
5 792 461 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
5.89948e-315 5.36716e-315
0
13 Logic Switch~
5 633 806 0 10 11
0 57 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-5 -27 9 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
5.89948e-315 5.3568e-315
0
13 Logic Switch~
5 630 736 0 10 11
0 58 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3178 0 0
2
5.89948e-315 5.34643e-315
0
13 Logic Switch~
5 638 675 0 10 11
0 60 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -16 7 -8
2 B3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
5.89948e-315 5.32571e-315
0
13 Logic Switch~
5 640 627 0 1 11
0 59
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3951 0 0
2
5.89948e-315 5.30499e-315
0
13 Logic Switch~
5 631 885 0 10 11
0 56 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
4 Cin2
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8885 0 0
2
5.89948e-315 5.26354e-315
0
13 Logic Switch~
5 771 504 0 1 11
0 67
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3780 0 0
2
5.89948e-315 0
0
13 Logic Switch~
5 62 1170 0 1 11
0 78
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9265 0 0
2
5.89948e-315 5.37752e-315
0
13 Logic Switch~
5 61 1130 0 10 11
0 79 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9442 0 0
2
5.89948e-315 5.36716e-315
0
13 Logic Switch~
5 56 955 0 10 11
0 84 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
5.89948e-315 5.37752e-315
0
13 Logic Switch~
5 55 915 0 10 11
0 85 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.89948e-315 5.36716e-315
0
13 Logic Switch~
5 67 747 0 10 11
0 91 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9281 0 0
2
5.89948e-315 5.37752e-315
0
13 Logic Switch~
5 66 707 0 10 11
0 92 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8464 0 0
2
5.89948e-315 5.36716e-315
0
13 Logic Switch~
5 57 489 0 1 11
0 98
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
5.89948e-315 5.30499e-315
0
13 Logic Switch~
5 58 529 0 10 11
0 97 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3171 0 0
2
5.89948e-315 5.26354e-315
0
13 Logic Switch~
5 62 625 0 1 11
0 71
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4139 0 0
2
5.89948e-315 0
0
8 2-In OR~
219 194 161 0 3 22
0 2 3 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
6435 0 0
2
44059.4 0
0
9 2-In AND~
219 131 99 0 3 22
0 6 7 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
5283 0 0
2
44059.4 0
0
9 2-In AND~
219 133 196 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
6874 0 0
2
44059.4 0
0
9 Inverter~
13 72 176 0 2 22
0 7 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
5305 0 0
2
44059.4 0
0
14 Logic Display~
6 598 129 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
44059.4 6
0
9 2-In XOR~
219 538 147 0 3 22
0 11 12 10
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
969 0 0
2
44059.4 5
0
14 Logic Display~
6 621 218 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
44059.4 4
0
9 2-In AND~
219 488 245 0 3 22
0 11 12 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3751 0 0
2
44059.4 3
0
8 2-In OR~
219 565 236 0 3 22
0 14 13 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4292 0 0
2
44059.4 2
0
9 2-In AND~
219 384 199 0 3 22
0 15 8 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6118 0 0
2
44059.4 1
0
9 2-In XOR~
219 415 138 0 3 22
0 15 8 11
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
34 0 0
2
44059.4 0
0
14 Logic Display~
6 1120 155 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s4
-6 -22 8 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
44059.4 14
0
14 Logic Display~
6 1174 168 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
44059.4 13
0
14 Logic Display~
6 1237 193 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
44059.4 12
0
14 Logic Display~
6 1290 212 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
44059.4 11
0
14 Logic Display~
6 1141 261 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
44059.4 10
0
6 74LS83
105 1027 187 0 14 29
0 26 27 28 29 25 24 23 22 21
20 19 18 17 16
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6748 0 0
2
44059.4 9
0
9 2-In XOR~
219 335 1362 0 3 22
0 33 32 30
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6901 0 0
2
44059.4 5
0
9 2-In AND~
219 334 1451 0 3 22
0 33 32 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
842 0 0
2
44059.4 4
0
14 Logic Display~
6 405 1344 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
44059.4 3
0
14 Logic Display~
6 401 1433 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
44059.4 2
0
9 Inverter~
13 707 1268 0 2 22
0 38 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
4720 0 0
2
5.89948e-315 0
0
9 Inverter~
13 720 1207 0 2 22
0 39 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
5551 0 0
2
5.89948e-315 0
0
9 Inverter~
13 717 1148 0 2 22
0 41 36
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
6986 0 0
2
5.89948e-315 0
0
9 Inverter~
13 717 1090 0 2 22
0 40 37
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
8745 0 0
2
5.89948e-315 0
0
6 74LS83
105 938 1062 0 14 29
0 48 49 50 51 37 36 35 34 47
46 45 44 43 42
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U13
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9592 0 0
2
5.89948e-315 5.43451e-315
0
14 Logic Display~
6 991 1015 0 1 2
10 42
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.89948e-315 5.43192e-315
0
14 Logic Display~
6 1201 1087 0 1 2
10 43
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89948e-315 5.42933e-315
0
14 Logic Display~
6 1148 1068 0 1 2
10 44
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
5.89948e-315 5.42414e-315
0
14 Logic Display~
6 1085 1043 0 1 2
10 45
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9466 0 0
2
5.89948e-315 5.41896e-315
0
14 Logic Display~
6 1040 1028 0 1 2
10 46
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s5
-6 -22 8 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3266 0 0
2
5.89948e-315 5.41378e-315
0
9 2-In XOR~
219 724 814 0 3 22
0 57 56 52
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
7693 0 0
2
5.89948e-315 0
0
9 2-In XOR~
219 722 744 0 3 22
0 58 56 53
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3723 0 0
2
5.89948e-315 0
0
9 2-In XOR~
219 719 685 0 3 22
0 60 56 54
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3440 0 0
2
5.89948e-315 0
0
9 2-In XOR~
219 719 636 0 3 22
0 59 56 55
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
6263 0 0
2
5.89948e-315 0
0
14 Logic Display~
6 1046 567 0 1 2
10 65
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s4
-6 -22 8 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4900 0 0
2
5.89948e-315 5.41896e-315
0
14 Logic Display~
6 1100 580 0 1 2
10 64
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8783 0 0
2
5.89948e-315 5.41378e-315
0
14 Logic Display~
6 1163 605 0 1 2
10 63
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3221 0 0
2
5.89948e-315 5.4086e-315
0
14 Logic Display~
6 1216 624 0 1 2
10 62
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3215 0 0
2
5.89948e-315 5.40342e-315
0
14 Logic Display~
6 1013 560 0 1 2
10 61
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
5.89948e-315 5.39824e-315
0
6 74LS83
105 953 599 0 14 29
0 66 67 68 69 55 54 53 52 56
65 64 63 62 61
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U10
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7121 0 0
2
5.89948e-315 5.39306e-315
0
14 Logic Display~
6 398 1227 0 1 2
10 72
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
5.89948e-315 0
0
14 Logic Display~
6 459 1138 0 1 2
10 73
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
5.89948e-315 5.3568e-315
0
9 2-In XOR~
219 293 1156 0 3 22
0 74 75 73
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
7804 0 0
2
5.89948e-315 5.34643e-315
0
9 2-In AND~
219 243 1254 0 3 22
0 74 75 76
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
5523 0 0
2
5.89948e-315 5.32571e-315
0
8 2-In OR~
219 320 1245 0 3 22
0 77 76 72
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3330 0 0
2
5.89948e-315 5.30499e-315
0
9 2-In AND~
219 139 1208 0 3 22
0 79 78 77
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3465 0 0
2
5.89948e-315 5.26354e-315
0
9 2-In XOR~
219 170 1147 0 3 22
0 79 78 74
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8396 0 0
2
5.89948e-315 0
0
14 Logic Display~
6 453 923 0 1 2
10 80
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.89948e-315 5.3568e-315
0
9 2-In XOR~
219 287 941 0 3 22
0 81 70 80
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7849 0 0
2
5.89948e-315 5.34643e-315
0
9 2-In AND~
219 237 1039 0 3 22
0 81 70 82
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
6343 0 0
2
5.89948e-315 5.32571e-315
0
8 2-In OR~
219 314 1030 0 3 22
0 83 82 75
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7376 0 0
2
5.89948e-315 5.30499e-315
0
9 2-In AND~
219 133 993 0 3 22
0 85 84 83
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9156 0 0
2
5.89948e-315 5.26354e-315
0
9 2-In XOR~
219 164 932 0 3 22
0 85 84 81
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5776 0 0
2
5.89948e-315 0
0
14 Logic Display~
6 464 715 0 1 2
10 86
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
5.89948e-315 5.3568e-315
0
9 2-In XOR~
219 298 733 0 3 22
0 87 88 86
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4459 0 0
2
5.89948e-315 5.34643e-315
0
9 2-In AND~
219 248 831 0 3 22
0 87 88 89
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3760 0 0
2
5.89948e-315 5.32571e-315
0
8 2-In OR~
219 325 822 0 3 22
0 90 89 70
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
754 0 0
2
5.89948e-315 5.30499e-315
0
9 2-In AND~
219 144 785 0 3 22
0 92 91 90
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9767 0 0
2
5.89948e-315 5.26354e-315
0
9 2-In XOR~
219 175 724 0 3 22
0 92 91 87
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7978 0 0
2
5.89948e-315 0
0
9 2-In XOR~
219 166 506 0 3 22
0 98 97 94
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3142 0 0
2
5.89948e-315 5.39306e-315
0
9 2-In AND~
219 135 567 0 3 22
0 98 97 96
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3284 0 0
2
5.89948e-315 5.38788e-315
0
8 2-In OR~
219 316 604 0 3 22
0 96 95 88
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
659 0 0
2
5.89948e-315 5.37752e-315
0
9 2-In AND~
219 239 613 0 3 22
0 94 71 95
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3800 0 0
2
5.89948e-315 5.36716e-315
0
9 2-In XOR~
219 289 515 0 3 22
0 94 71 93
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6792 0 0
2
5.89948e-315 5.34643e-315
0
14 Logic Display~
6 455 497 0 1 2
10 93
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
5.89948e-315 5.32571e-315
0
126
3 1 2 0 0 4224 0 45 44 0 0 3
152 99
152 152
181 152
3 2 3 0 0 8320 0 46 44 0 0 3
154 196
154 170
181 170
1 2 4 0 0 8320 0 1 46 0 0 3
87 217
87 205
109 205
2 1 5 0 0 8320 0 47 46 0 0 3
93 176
93 187
109 187
1 1 6 0 0 4224 0 2 45 0 0 2
96 90
107 90
1 2 7 0 0 4224 0 14 45 0 0 4
41 142
82 142
82 108
107 108
0 2 8 0 0 4096 0 0 54 17 0 4
340 161
378 161
378 147
399 147
1 1 7 0 0 0 0 14 47 0 0 3
41 142
41 176
57 176
3 1 9 0 0 4224 0 52 50 0 0 2
598 236
621 236
3 1 10 0 0 4224 0 49 48 0 0 2
571 147
598 147
0 1 11 0 0 4096 0 0 49 16 0 2
464 138
522 138
0 2 12 0 0 4096 0 0 49 15 0 3
423 257
423 156
522 156
3 2 13 0 0 4224 0 51 52 0 0 2
509 245
552 245
3 1 14 0 0 4224 0 53 52 0 0 4
405 199
522 199
522 227
552 227
1 2 12 0 0 4224 0 3 51 0 0 4
323 257
444 257
444 254
464 254
3 1 11 0 0 8320 0 54 51 0 0 3
448 138
464 138
464 236
3 2 8 0 0 4224 0 44 53 0 0 4
227 161
340 161
340 208
360 208
0 1 15 0 0 4224 0 0 53 19 0 3
353 121
353 190
360 190
1 1 15 0 0 0 0 4 54 0 0 4
318 121
365 121
365 129
399 129
14 1 16 0 0 8320 0 60 59 0 0 4
1059 232
1098 232
1098 279
1141 279
13 1 17 0 0 4224 0 60 58 0 0 4
1059 205
1210 205
1210 230
1290 230
12 1 18 0 0 4224 0 60 57 0 0 4
1059 196
1223 196
1223 211
1237 211
11 1 19 0 0 8320 0 60 56 0 0 3
1059 187
1059 186
1174 186
10 1 20 0 0 4224 0 60 55 0 0 3
1059 178
1120 178
1120 173
1 9 21 0 0 8320 0 12 60 0 0 4
961 373
990 373
990 232
995 232
1 8 22 0 0 8320 0 8 60 0 0 4
858 343
903 343
903 214
995 214
1 7 23 0 0 12416 0 9 60 0 0 4
854 296
895 296
895 205
995 205
1 6 24 0 0 12416 0 10 60 0 0 4
852 253
888 253
888 196
995 196
1 5 25 0 0 12416 0 11 60 0 0 4
872 215
878 215
878 187
995 187
1 1 26 0 0 12416 0 7 60 0 0 4
878 49
886 49
886 151
995 151
1 2 27 0 0 12416 0 13 60 0 0 4
857 92
874 92
874 160
995 160
1 3 28 0 0 12416 0 6 60 0 0 4
848 138
861 138
861 169
995 169
1 4 29 0 0 12416 0 5 60 0 0 4
847 179
862 179
862 178
995 178
3 1 30 0 0 4224 0 61 63 0 0 2
368 1362
405 1362
3 1 31 0 0 4224 0 62 64 0 0 2
355 1451
401 1451
0 2 32 0 0 4096 0 0 62 38 0 3
243 1371
243 1460
310 1460
0 1 33 0 0 4096 0 0 62 39 0 3
263 1353
263 1442
310 1442
1 2 32 0 0 12416 0 16 61 0 0 4
203 1403
217 1403
217 1371
319 1371
1 1 33 0 0 4224 0 15 61 0 0 2
203 1353
319 1353
2 8 34 0 0 8320 0 65 69 0 0 4
728 1268
810 1268
810 1089
906 1089
2 7 35 0 0 8320 0 66 69 0 0 4
741 1207
795 1207
795 1080
906 1080
2 6 36 0 0 12416 0 67 69 0 0 4
738 1148
781 1148
781 1071
906 1071
2 5 37 0 0 12416 0 68 69 0 0 4
738 1090
768 1090
768 1062
906 1062
1 1 38 0 0 8320 0 22 65 0 0 3
630 1269
630 1268
692 1268
1 1 39 0 0 8320 0 21 66 0 0 3
627 1199
627 1207
705 1207
1 1 40 0 0 4224 0 19 68 0 0 2
637 1090
702 1090
1 1 41 0 0 8320 0 20 67 0 0 3
635 1138
635 1148
702 1148
14 1 42 0 0 8320 0 69 70 0 0 4
970 1107
1009 1107
1009 1033
991 1033
13 1 43 0 0 4224 0 69 71 0 0 4
970 1080
1121 1080
1121 1105
1201 1105
12 1 44 0 0 4224 0 69 72 0 0 4
970 1071
1134 1071
1134 1086
1148 1086
11 1 45 0 0 8320 0 69 73 0 0 3
970 1062
970 1061
1085 1061
10 1 46 0 0 4224 0 69 74 0 0 3
970 1053
1040 1053
1040 1046
1 9 47 0 0 4224 0 18 69 0 0 4
628 1348
901 1348
901 1107
906 1107
1 1 48 0 0 12416 0 23 69 0 0 4
789 924
797 924
797 1026
906 1026
1 2 49 0 0 12416 0 17 69 0 0 4
768 967
785 967
785 1035
906 1035
1 3 50 0 0 12416 0 24 69 0 0 4
759 1013
772 1013
772 1044
906 1044
1 4 51 0 0 12416 0 25 69 0 0 4
758 1054
773 1054
773 1053
906 1053
3 8 52 0 0 8320 0 75 84 0 0 4
757 814
825 814
825 626
921 626
3 7 53 0 0 8320 0 76 84 0 0 4
755 744
810 744
810 617
921 617
3 6 54 0 0 12416 0 77 84 0 0 4
752 685
796 685
796 608
921 608
3 5 55 0 0 12416 0 78 84 0 0 4
752 636
783 636
783 599
921 599
0 2 56 0 0 8192 0 0 75 65 0 3
688 824
688 823
708 823
0 2 56 0 0 0 0 0 76 65 0 2
688 753
706 753
0 2 56 0 0 0 0 0 77 65 0 3
688 692
688 694
703 694
0 2 56 0 0 4096 0 0 78 75 0 3
688 885
688 645
703 645
1 1 57 0 0 8320 0 29 75 0 0 3
645 806
645 805
708 805
1 1 58 0 0 8320 0 30 76 0 0 3
642 736
642 735
706 735
1 1 59 0 0 4224 0 32 78 0 0 2
652 627
703 627
1 1 60 0 0 8320 0 31 77 0 0 3
650 675
650 676
703 676
14 1 61 0 0 8320 0 84 83 0 0 4
985 644
1024 644
1024 578
1013 578
13 1 62 0 0 4224 0 84 82 0 0 4
985 617
1136 617
1136 642
1216 642
12 1 63 0 0 4224 0 84 81 0 0 4
985 608
1149 608
1149 623
1163 623
11 1 64 0 0 8320 0 84 80 0 0 3
985 599
985 598
1100 598
10 1 65 0 0 4224 0 84 79 0 0 3
985 590
1046 590
1046 585
1 9 56 0 0 4224 0 33 84 0 0 4
643 885
916 885
916 644
921 644
1 1 66 0 0 12416 0 28 84 0 0 4
804 461
812 461
812 563
921 563
1 2 67 0 0 12416 0 34 84 0 0 4
783 504
800 504
800 572
921 572
1 3 68 0 0 12416 0 27 84 0 0 4
774 550
787 550
787 581
921 581
1 4 69 0 0 12416 0 26 84 0 0 4
773 591
788 591
788 590
921 590
2 0 70 0 0 8192 0 93 0 0 104 3
271 950
183 950
183 1048
0 2 71 0 0 12288 0 0 107 119 0 4
173 625
189 625
189 622
215 622
3 1 72 0 0 4224 0 0 85 83 0 2
375 1245
398 1245
3 0 72 0 0 0 0 89 0 0 82 2
353 1245
376 1245
3 1 73 0 0 4224 0 87 86 0 0 2
326 1156
459 1156
0 1 74 0 0 4096 0 0 87 90 0 2
219 1147
277 1147
0 2 75 0 0 8192 0 0 87 89 0 3
178 1263
178 1165
277 1165
3 2 76 0 0 4224 0 88 89 0 0 2
264 1254
307 1254
3 1 77 0 0 4224 0 90 89 0 0 4
160 1208
277 1208
277 1236
307 1236
3 2 75 0 0 12416 0 95 88 0 0 6
347 1030
370 1030
370 1093
33 1093
33 1263
219 1263
3 1 74 0 0 8320 0 91 88 0 0 3
203 1147
219 1147
219 1245
0 2 78 0 0 4224 0 0 90 93 0 3
95 1170
95 1217
115 1217
0 1 79 0 0 4224 0 0 90 94 0 3
108 1130
108 1199
115 1199
1 2 78 0 0 0 0 35 91 0 0 4
74 1170
120 1170
120 1156
154 1156
1 1 79 0 0 0 0 36 91 0 0 4
73 1130
120 1130
120 1138
154 1138
3 1 80 0 0 4224 0 93 92 0 0 2
320 941
453 941
0 1 81 0 0 4096 0 0 93 99 0 2
213 932
271 932
3 2 82 0 0 4224 0 94 95 0 0 2
258 1039
301 1039
3 1 83 0 0 4224 0 96 95 0 0 4
154 993
271 993
271 1021
301 1021
3 1 81 0 0 8320 0 97 94 0 0 3
197 932
213 932
213 1030
0 2 84 0 0 4224 0 0 96 102 0 3
89 955
89 1002
109 1002
0 1 85 0 0 4224 0 0 96 103 0 3
102 915
102 984
109 984
1 2 84 0 0 0 0 37 97 0 0 4
68 955
114 955
114 941
148 941
1 1 85 0 0 0 0 38 97 0 0 4
67 915
114 915
114 923
148 923
3 2 70 0 0 12416 0 101 94 0 0 6
358 822
381 822
381 881
34 881
34 1048
213 1048
3 1 86 0 0 4224 0 99 98 0 0 2
331 733
464 733
0 1 87 0 0 4096 0 0 99 111 0 2
224 724
282 724
0 2 88 0 0 8192 0 0 99 110 0 3
183 840
183 742
282 742
3 2 89 0 0 4224 0 100 101 0 0 2
269 831
312 831
3 1 90 0 0 4224 0 102 101 0 0 4
165 785
282 785
282 813
312 813
0 2 88 0 0 8320 0 0 100 0 0 5
372 607
372 671
37 671
37 840
224 840
3 1 87 0 0 8320 0 103 100 0 0 3
208 724
224 724
224 822
0 2 91 0 0 4224 0 0 102 114 0 3
100 747
100 794
120 794
0 1 92 0 0 4224 0 0 102 115 0 3
113 707
113 776
120 776
1 2 91 0 0 0 0 39 103 0 0 4
79 747
125 747
125 733
159 733
1 1 92 0 0 0 0 40 103 0 0 4
78 707
125 707
125 715
159 715
3 0 88 0 0 0 0 106 0 0 110 3
349 604
372 604
372 607
3 1 93 0 0 4224 0 108 109 0 0 2
322 515
455 515
0 1 94 0 0 4096 0 0 108 122 0 2
215 506
273 506
1 2 71 0 0 8320 0 43 108 0 0 4
74 625
174 625
174 524
273 524
3 2 95 0 0 4224 0 107 106 0 0 2
260 613
303 613
3 1 96 0 0 4224 0 105 106 0 0 4
156 567
273 567
273 595
303 595
3 1 94 0 0 8320 0 104 107 0 0 3
199 506
215 506
215 604
0 2 97 0 0 4224 0 0 105 125 0 3
91 529
91 576
111 576
0 1 98 0 0 4224 0 0 105 126 0 3
104 489
104 558
111 558
1 2 97 0 0 0 0 42 104 0 0 4
70 529
116 529
116 515
150 515
1 1 98 0 0 0 0 41 104 0 0 4
69 489
116 489
116 497
150 497
93
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
563 146 582 170
568 152 576 168
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
512 159 533 183
518 164 526 180
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
605 137 644 161
612 143 636 159
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
626 229 673 253
633 235 665 251
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
502 241 521 265
507 247 515 263
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
453 257 474 281
459 262 467 278
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
448 215 467 239
453 221 461 237
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
512 108 531 132
517 114 525 130
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
398 177 417 201
403 182 411 198
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
593 214 612 238
598 219 606 235
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
441 114 460 138
446 119 454 135
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
539 250 558 274
544 255 552 271
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
349 209 368 233
354 214 362 230
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
390 149 409 173
395 154 403 170
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
538 203 559 227
544 209 552 225
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
351 162 372 186
357 168 365 184
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
389 97 410 121
395 103 403 119
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1149 280 1196 304
1156 286 1188 302
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
305 1324 326 1348
311 1330 319 1346
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
306 1375 325 1399
311 1380 319 1396
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
360 1367 379 1391
365 1372 373 1388
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
301 1414 322 1438
307 1420 315 1436
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
302 1463 321 1487
307 1468 315 1484
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
349 1427 368 1451
354 1432 362 1448
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
413 1351 452 1375
420 1356 444 1372
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
407 1443 462 1467
414 1449 454 1465
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
140 465 161 489
146 471 154 487
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
102 530 123 554
108 536 116 552
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
289 571 310 595
295 577 303 593
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
141 517 160 541
146 522 154 538
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
100 577 119 601
105 582 113 598
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
290 618 309 642
295 623 303 639
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
192 482 211 506
197 487 205 503
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
344 582 363 606
349 587 357 603
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
149 545 168 569
154 550 162 566
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
263 476 282 500
268 482 276 498
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
199 583 218 607
204 589 212 605
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
204 625 225 649
210 630 218 646
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
253 609 272 633
258 615 266 631
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
263 527 284 551
269 532 277 548
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
314 514 333 538
319 520 327 536
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
463 521 494 545
470 527 486 543
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
312 940 331 964
317 946 325 962
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
261 953 282 977
267 958 275 974
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
251 1035 270 1059
256 1041 264 1057
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
202 1051 223 1075
208 1056 216 1072
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
197 1009 216 1033
202 1015 210 1031
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
261 902 280 926
266 908 274 924
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
147 971 166 995
152 976 160 992
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
190 908 209 932
195 913 203 929
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
98 1003 117 1027
103 1008 111 1024
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
139 943 158 967
144 948 152 964
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
100 956 121 980
106 962 114 978
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
138 891 159 915
144 897 152 913
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
472 739 503 783
479 745 495 777
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
461 947 492 971
468 953 484 969
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
467 1162 498 1186
474 1167 490 1183
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
407 1238 454 1262
414 1244 446 1260
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
150 735 169 759
155 741 163 757
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
267 745 296 769
273 751 289 767
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
107 748 134 772
112 753 128 769
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
107 795 126 819
112 800 120 816
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
158 763 177 787
163 769 171 785
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
205 803 232 827
210 808 226 824
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
209 844 236 868
214 849 230 865
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
259 830 286 854
264 835 280 851
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
295 790 316 814
301 795 309 811
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
297 837 318 861
303 843 311 859
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
353 800 372 824
358 805 366 821
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
284 997 311 1021
289 1003 305 1019
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
288 1044 307 1068
293 1049 301 1065
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
342 1008 361 1032
347 1013 355 1029
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
290 1212 317 1236
295 1217 311 1233
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
291 1259 320 1283
297 1265 313 1281
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
345 1223 372 1247
350 1229 366 1245
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
145 1158 166 1182
151 1163 159 1179
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
265 694 296 718
272 699 288 715
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
319 732 350 756
326 737 342 753
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
147 683 174 707
152 689 168 705
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
198 699 221 723
205 705 213 721
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
141 1105 170 1129
147 1111 163 1127
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
193 1125 216 1149
200 1131 208 1147
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
263 1118 292 1142
269 1123 285 1139
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
263 1168 290 1192
268 1173 284 1189
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
315 1155 344 1179
321 1161 337 1177
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
104 1171 131 1195
109 1177 125 1193
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
104 1218 123 1242
109 1223 117 1239
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
153 1186 174 1210
159 1191 167 1207
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
198 1228 225 1252
203 1233 219 1249
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
208 1266 235 1290
213 1271 229 1287
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
253 1250 280 1274
258 1255 274 1271
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
989 513 1036 537
996 519 1028 535
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1055 1160 1102 1184
1062 1166 1094 1182
4 Cout
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
