CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
550 490 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
103
13 Logic Switch~
5 756 967 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44038.4 8
0
13 Logic Switch~
5 616 1348 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
4 Cin3
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
44038.4 7
0
13 Logic Switch~
5 625 1090 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44038.4 6
0
13 Logic Switch~
5 623 1138 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -16 7 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
44038.4 5
0
13 Logic Switch~
5 615 1199 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
44038.4 4
0
13 Logic Switch~
5 618 1269 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-5 -30 9 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
44038.4 3
0
13 Logic Switch~
5 777 924 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
44038.4 2
0
13 Logic Switch~
5 747 1013 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
44038.4 1
0
13 Logic Switch~
5 746 1054 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
44038.4 0
0
13 Logic Switch~
5 761 591 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
44038.4 8
0
13 Logic Switch~
5 762 550 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
44038.4 7
0
13 Logic Switch~
5 792 461 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
44038.4 6
0
13 Logic Switch~
5 633 806 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-5 -27 9 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
44038.4 5
0
13 Logic Switch~
5 630 736 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
44038.4 4
0
13 Logic Switch~
5 638 675 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -16 7 -8
2 B3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
44038.4 3
0
13 Logic Switch~
5 640 627 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
44038.4 2
0
13 Logic Switch~
5 631 885 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
4 Cin2
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5616 0 0
2
44038.4 1
0
13 Logic Switch~
5 771 504 0 1 11
0 35
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A3
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
44038.4 0
0
13 Logic Switch~
5 62 1170 0 1 11
0 46
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
44038.4 7
0
13 Logic Switch~
5 61 1130 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3108 0 0
2
44038.4 6
0
13 Logic Switch~
5 56 955 0 10 11
0 52 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4299 0 0
2
44038.4 7
0
13 Logic Switch~
5 55 915 0 10 11
0 53 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9672 0 0
2
44038.4 6
0
13 Logic Switch~
5 67 747 0 10 11
0 59 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7876 0 0
2
44038.4 7
0
13 Logic Switch~
5 66 707 0 10 11
0 60 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
44038.4 6
0
13 Logic Switch~
5 57 489 0 1 11
0 66
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
44038.4 2
0
13 Logic Switch~
5 58 529 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
44038.4 1
0
13 Logic Switch~
5 62 625 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
44038.4 0
0
13 Logic Switch~
5 646 109 0 10 11
0 78 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-5 -26 9 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 750 390 0 1 11
0 72
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 Cin1
-12 -26 16 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
961 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 661 232 0 1 11
0 76
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 641 270 0 10 11
0 75 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 643 313 0 10 11
0 74 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3951 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 647 360 0 1 11
0 73
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 B1
-5 -27 9 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 667 66 0 10 11
0 77 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3780 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 637 155 0 1 11
0 79
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9265 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 636 196 0 1 11
0 80
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 63 399 0 10 11
0 84 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 59 303 0 1 11
0 87
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 58 263 0 1 11
0 88
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 51 136 0 1 11
0 91
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8464 0 0
2
5.89947e-315 0
0
13 Logic Switch~
5 51 86 0 10 11
0 92 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7168 0 0
2
5.89947e-315 0
0
9 Inverter~
13 707 1268 0 2 22
0 6 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
3171 0 0
2
44038.4 0
0
9 Inverter~
13 720 1207 0 2 22
0 7 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 10 0
1 U
4139 0 0
2
44038.4 0
0
9 Inverter~
13 717 1148 0 2 22
0 9 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 10 0
1 U
6435 0 0
2
44038.4 0
0
9 Inverter~
13 717 1090 0 2 22
0 8 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U12A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
5283 0 0
2
44038.4 0
0
6 74LS83
105 938 1062 0 14 29
0 16 17 18 19 5 4 3 2 15
14 13 12 11 10
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U13
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6874 0 0
2
44038.4 18
0
14 Logic Display~
6 991 1015 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
44038.4 17
0
14 Logic Display~
6 1201 1087 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
44038.4 16
0
14 Logic Display~
6 1148 1068 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
44038.4 15
0
14 Logic Display~
6 1085 1043 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
44038.4 14
0
14 Logic Display~
6 1040 1028 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s5
-6 -22 8 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
44038.4 13
0
9 2-In XOR~
219 724 814 0 3 22
0 25 24 20
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
4292 0 0
2
44038.4 0
0
9 2-In XOR~
219 722 744 0 3 22
0 26 24 21
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
6118 0 0
2
44038.4 0
0
9 2-In XOR~
219 719 685 0 3 22
0 28 24 22
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
34 0 0
2
44038.4 0
0
9 2-In XOR~
219 719 636 0 3 22
0 27 24 23
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
6357 0 0
2
44038.4 0
0
14 Logic Display~
6 1046 567 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s4
-6 -22 8 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
44038.4 14
0
14 Logic Display~
6 1100 580 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
44038.4 13
0
14 Logic Display~
6 1163 605 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
44038.4 12
0
14 Logic Display~
6 1216 624 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
44038.4 11
0
14 Logic Display~
6 1013 560 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
44038.4 10
0
6 74LS83
105 953 599 0 14 29
0 34 35 36 37 23 22 21 20 24
33 32 31 30 29
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U10
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6901 0 0
2
44038.4 9
0
14 Logic Display~
6 398 1227 0 1 2
10 40
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
44038.4 0
0
14 Logic Display~
6 459 1138 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
44038.4 5
0
9 2-In XOR~
219 293 1156 0 3 22
0 42 43 41
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
4212 0 0
2
44038.4 4
0
9 2-In AND~
219 243 1254 0 3 22
0 42 43 44
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
4720 0 0
2
44038.4 3
0
8 2-In OR~
219 320 1245 0 3 22
0 45 44 40
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
5551 0 0
2
44038.4 2
0
9 2-In AND~
219 139 1208 0 3 22
0 47 46 45
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6986 0 0
2
44038.4 1
0
9 2-In XOR~
219 170 1147 0 3 22
0 47 46 42
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8745 0 0
2
44038.4 0
0
14 Logic Display~
6 453 923 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
44038.4 5
0
9 2-In XOR~
219 287 941 0 3 22
0 49 38 48
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8748 0 0
2
44038.4 4
0
9 2-In AND~
219 237 1039 0 3 22
0 49 38 50
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7168 0 0
2
44038.4 3
0
8 2-In OR~
219 314 1030 0 3 22
0 51 50 43
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
631 0 0
2
44038.4 2
0
9 2-In AND~
219 133 993 0 3 22
0 53 52 51
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9466 0 0
2
44038.4 1
0
9 2-In XOR~
219 164 932 0 3 22
0 53 52 49
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3266 0 0
2
44038.4 0
0
14 Logic Display~
6 464 715 0 1 2
10 54
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
44038.4 5
0
9 2-In XOR~
219 298 733 0 3 22
0 55 56 54
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3723 0 0
2
44038.4 4
0
9 2-In AND~
219 248 831 0 3 22
0 55 56 57
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3440 0 0
2
44038.4 3
0
8 2-In OR~
219 325 822 0 3 22
0 58 57 38
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6263 0 0
2
44038.4 2
0
9 2-In AND~
219 144 785 0 3 22
0 60 59 58
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4900 0 0
2
44038.4 1
0
9 2-In XOR~
219 175 724 0 3 22
0 60 59 55
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8783 0 0
2
44038.4 0
0
9 2-In XOR~
219 166 506 0 3 22
0 66 65 62
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3221 0 0
2
44038.4 9
0
9 2-In AND~
219 135 567 0 3 22
0 66 65 64
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3215 0 0
2
44038.4 8
0
8 2-In OR~
219 316 604 0 3 22
0 64 63 56
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7903 0 0
2
44038.4 7
0
9 2-In AND~
219 239 613 0 3 22
0 62 39 63
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7121 0 0
2
44038.4 6
0
9 2-In XOR~
219 289 515 0 3 22
0 62 39 61
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4484 0 0
2
44038.4 4
0
14 Logic Display~
6 455 497 0 1 2
10 61
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
44038.4 3
0
6 74LS83
105 828 204 0 14 29
0 77 78 79 80 76 75 74 73 72
71 70 69 68 67
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7804 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 942 278 0 1 2
10 67
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 1091 229 0 1 2
10 68
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 1038 210 0 1 2
10 69
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 975 185 0 1 2
10 70
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 921 172 0 1 2
10 71
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 s4
-6 -22 8 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 350 271 0 1 2
10 82
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
5.89947e-315 0
0
9 2-In XOR~
219 290 289 0 3 22
0 83 84 82
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6343 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 373 360 0 1 2
10 81
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
5.89947e-315 0
0
9 2-In AND~
219 240 387 0 3 22
0 83 84 85
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9156 0 0
2
5.89947e-315 0
0
8 2-In OR~
219 317 378 0 3 22
0 86 85 81
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5776 0 0
2
5.89947e-315 0
0
9 2-In AND~
219 136 341 0 3 22
0 88 87 86
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7207 0 0
2
5.89947e-315 0
0
9 2-In XOR~
219 167 280 0 3 22
0 88 87 83
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4459 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 261 166 0 1 2
10 90
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
5.89947e-315 0
0
14 Logic Display~
6 265 77 0 1 2
10 89
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
5.89947e-315 0
0
9 2-In AND~
219 194 184 0 3 22
0 92 91 90
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9767 0 0
2
5.89947e-315 0
0
9 2-In XOR~
219 195 95 0 3 22
0 92 91 89
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7978 0 0
2
5.89947e-315 0
0
119
2 8 2 0 0 8336 0 42 46 0 0 4
728 1268
810 1268
810 1089
906 1089
2 7 3 0 0 8320 0 43 46 0 0 4
741 1207
795 1207
795 1080
906 1080
2 6 4 0 0 12416 0 44 46 0 0 4
738 1148
781 1148
781 1071
906 1071
2 5 5 0 0 12416 0 45 46 0 0 4
738 1090
768 1090
768 1062
906 1062
1 1 6 0 0 8320 0 6 42 0 0 3
630 1269
630 1268
692 1268
1 1 7 0 0 8320 0 5 43 0 0 3
627 1199
627 1207
705 1207
1 1 8 0 0 4224 0 3 45 0 0 2
637 1090
702 1090
1 1 9 0 0 8320 0 4 44 0 0 3
635 1138
635 1148
702 1148
14 1 10 0 0 8320 0 46 47 0 0 4
970 1107
1009 1107
1009 1033
991 1033
13 1 11 0 0 4224 0 46 48 0 0 4
970 1080
1121 1080
1121 1105
1201 1105
12 1 12 0 0 4224 0 46 49 0 0 4
970 1071
1134 1071
1134 1086
1148 1086
11 1 13 0 0 8320 0 46 50 0 0 3
970 1062
970 1061
1085 1061
10 1 14 0 0 4224 0 46 51 0 0 3
970 1053
1040 1053
1040 1046
1 9 15 0 0 4224 0 2 46 0 0 4
628 1348
901 1348
901 1107
906 1107
1 1 16 0 0 12416 0 7 46 0 0 4
789 924
797 924
797 1026
906 1026
1 2 17 0 0 12416 0 1 46 0 0 4
768 967
785 967
785 1035
906 1035
1 3 18 0 0 12416 0 8 46 0 0 4
759 1013
772 1013
772 1044
906 1044
1 4 19 0 0 12416 0 9 46 0 0 4
758 1054
773 1054
773 1053
906 1053
3 8 20 0 0 8320 0 52 61 0 0 4
757 814
825 814
825 626
921 626
3 7 21 0 0 8320 0 53 61 0 0 4
755 744
810 744
810 617
921 617
3 6 22 0 0 12416 0 54 61 0 0 4
752 685
796 685
796 608
921 608
3 5 23 0 0 12416 0 55 61 0 0 4
752 636
783 636
783 599
921 599
0 2 24 0 0 8192 0 0 52 26 0 3
688 824
688 823
708 823
0 2 24 0 0 0 0 0 53 26 0 2
688 753
706 753
0 2 24 0 0 0 0 0 54 26 0 3
688 692
688 694
703 694
0 2 24 0 0 4096 0 0 55 36 0 3
688 885
688 645
703 645
1 1 25 0 0 8320 0 13 52 0 0 3
645 806
645 805
708 805
1 1 26 0 0 8320 0 14 53 0 0 3
642 736
642 735
706 735
1 1 27 0 0 4224 0 16 55 0 0 2
652 627
703 627
1 1 28 0 0 8320 0 15 54 0 0 3
650 675
650 676
703 676
14 1 29 0 0 8320 0 61 60 0 0 4
985 644
1024 644
1024 578
1013 578
13 1 30 0 0 4224 0 61 59 0 0 4
985 617
1136 617
1136 642
1216 642
12 1 31 0 0 4224 0 61 58 0 0 4
985 608
1149 608
1149 623
1163 623
11 1 32 0 0 8320 0 61 57 0 0 3
985 599
985 598
1100 598
10 1 33 0 0 4224 0 61 56 0 0 3
985 590
1046 590
1046 585
1 9 24 0 0 4224 0 17 61 0 0 4
643 885
916 885
916 644
921 644
1 1 34 0 0 12416 0 12 61 0 0 4
804 461
812 461
812 563
921 563
1 2 35 0 0 12416 0 18 61 0 0 4
783 504
800 504
800 572
921 572
1 3 36 0 0 12416 0 11 61 0 0 4
774 550
787 550
787 581
921 581
1 4 37 0 0 12416 0 10 61 0 0 4
773 591
788 591
788 590
921 590
2 0 38 0 0 8192 0 70 0 0 65 3
271 950
183 950
183 1048
0 2 39 0 0 12288 0 0 84 80 0 4
173 625
189 625
189 622
215 622
3 1 40 0 0 4224 0 0 62 44 0 2
375 1245
398 1245
3 0 40 0 0 0 0 66 0 0 43 2
353 1245
376 1245
3 1 41 0 0 4224 0 64 63 0 0 2
326 1156
459 1156
0 1 42 0 0 4096 0 0 64 51 0 2
219 1147
277 1147
0 2 43 0 0 8192 0 0 64 50 0 3
178 1263
178 1165
277 1165
3 2 44 0 0 4224 0 65 66 0 0 2
264 1254
307 1254
3 1 45 0 0 4224 0 67 66 0 0 4
160 1208
277 1208
277 1236
307 1236
3 2 43 0 0 12416 0 72 65 0 0 6
347 1030
370 1030
370 1093
33 1093
33 1263
219 1263
3 1 42 0 0 8320 0 68 65 0 0 3
203 1147
219 1147
219 1245
0 2 46 0 0 4224 0 0 67 54 0 3
95 1170
95 1217
115 1217
0 1 47 0 0 4224 0 0 67 55 0 3
108 1130
108 1199
115 1199
1 2 46 0 0 0 0 19 68 0 0 4
74 1170
120 1170
120 1156
154 1156
1 1 47 0 0 0 0 20 68 0 0 4
73 1130
120 1130
120 1138
154 1138
3 1 48 0 0 4224 0 70 69 0 0 2
320 941
453 941
0 1 49 0 0 4096 0 0 70 60 0 2
213 932
271 932
3 2 50 0 0 4224 0 71 72 0 0 2
258 1039
301 1039
3 1 51 0 0 4224 0 73 72 0 0 4
154 993
271 993
271 1021
301 1021
3 1 49 0 0 8320 0 74 71 0 0 3
197 932
213 932
213 1030
0 2 52 0 0 4224 0 0 73 63 0 3
89 955
89 1002
109 1002
0 1 53 0 0 4224 0 0 73 64 0 3
102 915
102 984
109 984
1 2 52 0 0 0 0 21 74 0 0 4
68 955
114 955
114 941
148 941
1 1 53 0 0 0 0 22 74 0 0 4
67 915
114 915
114 923
148 923
3 2 38 0 0 12416 0 78 71 0 0 6
358 822
381 822
381 881
34 881
34 1048
213 1048
3 1 54 0 0 4224 0 76 75 0 0 2
331 733
464 733
0 1 55 0 0 4096 0 0 76 72 0 2
224 724
282 724
0 2 56 0 0 8192 0 0 76 71 0 3
183 840
183 742
282 742
3 2 57 0 0 4224 0 77 78 0 0 2
269 831
312 831
3 1 58 0 0 4224 0 79 78 0 0 4
165 785
282 785
282 813
312 813
0 2 56 0 0 8320 0 0 77 0 0 5
372 607
372 671
37 671
37 840
224 840
3 1 55 0 0 8320 0 80 77 0 0 3
208 724
224 724
224 822
0 2 59 0 0 4224 0 0 79 75 0 3
100 747
100 794
120 794
0 1 60 0 0 4224 0 0 79 76 0 3
113 707
113 776
120 776
1 2 59 0 0 0 0 23 80 0 0 4
79 747
125 747
125 733
159 733
1 1 60 0 0 0 0 24 80 0 0 4
78 707
125 707
125 715
159 715
3 0 56 0 0 0 0 83 0 0 71 3
349 604
372 604
372 607
3 1 61 0 0 4224 0 85 86 0 0 2
322 515
455 515
0 1 62 0 0 4096 0 0 85 83 0 2
215 506
273 506
1 2 39 0 0 8320 0 27 85 0 0 4
74 625
174 625
174 524
273 524
3 2 63 0 0 4224 0 84 83 0 0 2
260 613
303 613
3 1 64 0 0 4224 0 82 83 0 0 4
156 567
273 567
273 595
303 595
3 1 62 0 0 8320 0 81 84 0 0 3
199 506
215 506
215 604
0 2 65 0 0 4224 0 0 82 86 0 3
91 529
91 576
111 576
0 1 66 0 0 4224 0 0 82 87 0 3
104 489
104 558
111 558
1 2 65 0 0 0 0 26 81 0 0 4
70 529
116 529
116 515
150 515
1 1 66 0 0 0 0 25 81 0 0 4
69 489
116 489
116 497
150 497
14 1 67 0 0 8320 0 87 88 0 0 4
860 249
899 249
899 296
942 296
13 1 68 0 0 4224 0 87 89 0 0 4
860 222
1011 222
1011 247
1091 247
12 1 69 0 0 4224 0 87 90 0 0 4
860 213
1024 213
1024 228
1038 228
11 1 70 0 0 8320 0 87 91 0 0 3
860 204
860 203
975 203
10 1 71 0 0 4224 0 87 92 0 0 3
860 195
921 195
921 190
1 9 72 0 0 8320 0 29 87 0 0 4
762 390
791 390
791 249
796 249
1 8 73 0 0 8320 0 33 87 0 0 4
659 360
704 360
704 231
796 231
1 7 74 0 0 12416 0 32 87 0 0 4
655 313
696 313
696 222
796 222
1 6 75 0 0 12416 0 31 87 0 0 4
653 270
689 270
689 213
796 213
1 5 76 0 0 12416 0 30 87 0 0 4
673 232
679 232
679 204
796 204
1 1 77 0 0 12416 0 34 87 0 0 4
679 66
687 66
687 168
796 168
1 2 78 0 0 12416 0 28 87 0 0 4
658 109
675 109
675 177
796 177
1 3 79 0 0 12416 0 35 87 0 0 4
649 155
662 155
662 186
796 186
1 4 80 0 0 12416 0 36 87 0 0 4
648 196
663 196
663 195
796 195
3 1 81 0 0 4224 0 97 95 0 0 2
350 378
373 378
3 1 82 0 0 4224 0 94 93 0 0 2
323 289
350 289
0 1 83 0 0 4096 0 0 94 109 0 2
216 280
274 280
0 2 84 0 0 4096 0 0 94 108 0 3
175 399
175 298
274 298
3 2 85 0 0 4224 0 96 97 0 0 2
261 387
304 387
3 1 86 0 0 4224 0 98 97 0 0 4
157 341
274 341
274 369
304 369
1 2 84 0 0 4224 0 37 96 0 0 4
75 399
196 399
196 396
216 396
3 1 83 0 0 8320 0 99 96 0 0 3
200 280
216 280
216 378
0 2 87 0 0 4224 0 0 98 112 0 3
92 303
92 350
112 350
0 1 88 0 0 4224 0 0 98 113 0 3
105 263
105 332
112 332
1 2 87 0 0 0 0 38 99 0 0 4
71 303
117 303
117 289
151 289
1 1 88 0 0 0 0 39 99 0 0 4
70 263
117 263
117 271
151 271
3 1 89 0 0 4224 0 103 101 0 0 2
228 95
265 95
3 1 90 0 0 4224 0 102 100 0 0 2
215 184
261 184
0 2 91 0 0 4096 0 0 102 118 0 3
103 104
103 193
170 193
0 1 92 0 0 4096 0 0 102 119 0 3
123 86
123 175
170 175
1 2 91 0 0 12416 0 40 103 0 0 4
63 136
77 136
77 104
179 104
1 1 92 0 0 4224 0 41 103 0 0 2
63 86
179 86
93
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1055 1160 1102 1184
1062 1166 1094 1182
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1070 697 1117 721
1077 703 1109 719
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
950 297 997 321
957 303 989 319
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
253 1250 280 1274
258 1255 274 1271
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
208 1266 235 1290
213 1271 229 1287
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
198 1228 225 1252
203 1233 219 1249
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
153 1186 174 1210
159 1191 167 1207
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
104 1218 123 1242
109 1223 117 1239
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
104 1171 131 1195
109 1177 125 1193
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
315 1155 344 1179
321 1161 337 1177
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
263 1168 290 1192
268 1173 284 1189
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
263 1118 292 1142
269 1123 285 1139
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
193 1125 216 1149
200 1131 208 1147
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
141 1105 170 1129
147 1111 163 1127
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
198 699 221 723
205 705 213 721
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
147 683 174 707
152 689 168 705
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
319 732 350 756
326 737 342 753
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
265 694 296 718
272 699 288 715
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
145 1158 166 1182
151 1163 159 1179
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
345 1223 372 1247
350 1229 366 1245
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
291 1259 320 1283
297 1265 313 1281
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
290 1212 317 1236
295 1217 311 1233
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
342 1008 361 1032
347 1013 355 1029
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
288 1044 307 1068
293 1049 301 1065
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
284 997 311 1021
289 1003 305 1019
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
353 800 372 824
358 805 366 821
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
297 837 318 861
303 843 311 859
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
295 790 316 814
301 795 309 811
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
259 830 286 854
264 835 280 851
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
209 844 236 868
214 849 230 865
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
205 803 232 827
210 808 226 824
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
158 763 177 787
163 769 171 785
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
107 795 126 819
112 800 120 816
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
107 748 134 772
112 753 128 769
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
267 745 296 769
273 751 289 767
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
150 735 169 759
155 741 163 757
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
407 1238 454 1262
414 1244 446 1260
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
467 1162 498 1186
474 1167 490 1183
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
461 947 492 971
468 953 484 969
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
472 739 503 783
479 745 495 777
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
138 891 159 915
144 897 152 913
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
100 956 121 980
106 962 114 978
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
139 943 158 967
144 948 152 964
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
98 1003 117 1027
103 1008 111 1024
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
190 908 209 932
195 913 203 929
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
147 971 166 995
152 976 160 992
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
261 902 280 926
266 908 274 924
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
197 1009 216 1033
202 1015 210 1031
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
202 1051 223 1075
208 1056 216 1072
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
251 1035 270 1059
256 1041 264 1057
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
261 953 282 977
267 958 275 974
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
312 940 331 964
317 946 325 962
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
463 521 494 545
470 527 486 543
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
314 514 333 538
319 520 327 536
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
263 527 284 551
269 532 277 548
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
253 609 272 633
258 615 266 631
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
204 625 225 649
210 630 218 646
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
199 583 218 607
204 589 212 605
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
263 476 282 500
268 482 276 498
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
149 545 168 569
154 550 162 566
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
344 582 363 606
349 587 357 603
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
192 482 211 506
197 487 205 503
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
290 618 309 642
295 623 303 639
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
100 577 119 601
105 582 113 598
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
141 517 160 541
146 522 154 538
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
289 571 310 595
295 577 303 593
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
102 530 123 554
108 536 116 552
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
140 465 161 489
146 471 154 487
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
141 239 162 263
147 245 155 261
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
103 304 124 328
109 310 117 326
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
290 345 311 369
296 351 304 367
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
165 57 186 81
171 63 179 79
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
166 108 185 132
171 113 179 129
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
142 291 161 315
147 296 155 312
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
101 351 120 375
106 356 114 372
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
291 392 310 416
296 397 304 413
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
220 100 239 124
225 105 233 121
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
193 256 212 280
198 261 206 277
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
345 356 364 380
350 361 358 377
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
150 319 169 343
155 324 163 340
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
264 250 283 274
269 256 277 272
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
200 357 219 381
205 363 213 379
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
161 147 182 171
167 153 175 169
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
162 196 181 220
167 201 175 217
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
209 160 228 184
214 165 222 181
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
205 399 226 423
211 404 219 420
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
254 383 273 407
259 389 267 405
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
382 371 429 395
389 377 421 393
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
357 279 396 303
364 285 388 301
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
273 84 312 108
280 89 304 105
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
267 176 322 200
274 182 314 198
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
264 301 285 325
270 306 278 322
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
315 288 334 312
320 294 328 310
1 6
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
