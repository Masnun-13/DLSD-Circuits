CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 375 357 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 375 315 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 375 240 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3951 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 374 147 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 372 80 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3780 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 48 379 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9265 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 48 287 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 46 219 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9424 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 45 184 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.89946e-315 0
0
13 Logic Switch~
5 46 84 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
5.89946e-315 0
0
14 Logic Display~
6 616 315 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.89946e-315 0
0
9 2-In NOR~
219 542 333 0 3 22
0 3 3 2
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7168 0 0
2
5.89946e-315 0
0
9 2-In NOR~
219 444 324 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3171 0 0
2
5.89946e-315 0
0
14 Logic Display~
6 618 171 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.89946e-315 0
0
9 2-In NOR~
219 536 189 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
6435 0 0
2
5.89946e-315 0
0
9 2-In NOR~
219 442 231 0 3 22
0 9 9 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
5283 0 0
2
5.89946e-315 0
0
9 2-In NOR~
219 438 156 0 3 22
0 10 10 8
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6874 0 0
2
5.89946e-315 5.26354e-315
0
14 Logic Display~
6 512 71 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.89946e-315 0
0
9 2-In NOR~
219 436 89 0 3 22
0 12 12 11
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
34 0 0
2
5.89946e-315 0
0
14 Logic Display~
6 277 309 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.89946e-315 0
0
10 2-In NAND~
219 209 327 0 3 22
0 15 14 13
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8402 0 0
2
5.89946e-315 0
0
10 2-In NAND~
219 112 370 0 3 22
0 16 16 14
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3751 0 0
2
5.89946e-315 0
0
10 2-In NAND~
219 109 296 0 3 22
0 17 17 15
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4292 0 0
2
5.89946e-315 0
0
14 Logic Display~
6 269 189 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.89946e-315 0
0
10 2-In NAND~
219 212 207 0 3 22
0 19 19 18
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
34 0 0
2
5.89946e-315 0
0
10 2-In NAND~
219 124 198 0 3 22
0 21 20 19
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6357 0 0
2
5.89946e-315 0
0
14 Logic Display~
6 182 75 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
5.89946e-315 0
0
10 2-In NAND~
219 137 93 0 3 22
0 23 23 22
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3976 0 0
2
5.89946e-315 0
0
30
3 1 2 0 0 4224 0 12 11 0 0 2
581 333
616 333
0 2 3 0 0 8192 0 0 12 3 0 3
497 324
497 342
529 342
3 1 3 0 0 4224 0 13 12 0 0 2
483 324
529 324
1 2 4 0 0 12416 0 1 13 0 0 4
387 357
404 357
404 333
431 333
1 1 5 0 0 4224 0 2 13 0 0 2
387 315
431 315
3 1 6 0 0 4224 0 15 14 0 0 2
575 189
618 189
3 2 7 0 0 8320 0 16 15 0 0 4
481 231
507 231
507 198
523 198
3 1 8 0 0 4224 0 17 15 0 0 4
477 156
507 156
507 180
523 180
0 1 9 0 0 8192 0 0 16 10 0 3
405 240
405 222
429 222
1 2 9 0 0 4224 0 3 16 0 0 2
387 240
429 240
0 2 10 0 0 8192 0 0 17 12 0 3
403 147
403 165
425 165
1 1 10 0 0 4224 0 4 17 0 0 2
386 147
425 147
3 1 11 0 0 4224 0 19 18 0 0 2
475 89
512 89
0 2 12 0 0 8192 0 0 19 15 0 3
401 80
401 98
423 98
1 1 12 0 0 4224 0 5 19 0 0 2
384 80
423 80
3 1 13 0 0 4224 0 21 20 0 0 2
236 327
277 327
3 2 14 0 0 8320 0 22 21 0 0 4
139 370
163 370
163 336
185 336
3 1 15 0 0 4224 0 23 21 0 0 4
136 296
175 296
175 318
185 318
0 1 16 0 0 4096 0 0 22 20 0 3
75 379
75 361
88 361
1 2 16 0 0 4224 0 6 22 0 0 2
60 379
88 379
0 2 17 0 0 4096 0 0 23 22 0 3
71 287
71 305
85 305
1 1 17 0 0 4224 0 7 23 0 0 2
60 287
85 287
3 1 18 0 0 4224 0 25 24 0 0 2
239 207
269 207
0 1 19 0 0 4096 0 0 25 25 0 2
171 198
188 198
3 2 19 0 0 4224 0 26 25 0 0 4
151 198
171 198
171 216
188 216
1 2 20 0 0 4224 0 8 26 0 0 4
58 219
79 219
79 207
100 207
1 1 21 0 0 4224 0 9 26 0 0 4
57 184
79 184
79 189
100 189
3 1 22 0 0 4224 0 28 27 0 0 2
164 93
182 93
0 1 23 0 0 4096 0 0 28 30 0 2
89 84
113 84
1 2 23 0 0 4224 0 10 28 0 0 4
58 84
89 84
89 102
113 102
48
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
558 199 585 223
563 204 579 220
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
515 201 536 225
521 207 529 223
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
516 147 537 191
522 153 530 185
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
569 334 590 358
575 339 583 355
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 347 544 371
529 353 537 369
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
522 294 541 318
527 299 535 315
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
468 234 487 258
473 239 481 255
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
420 242 439 266
425 247 433 263
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
417 197 438 221
423 203 431 219
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
470 326 493 350
477 331 485 347
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
422 337 445 361
429 343 437 359
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
420 285 439 309
425 291 433 307
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
466 156 489 180
473 161 481 177
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
415 169 436 193
421 175 429 191
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
411 121 432 145
417 127 425 143
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
462 86 485 110
469 91 477 107
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
415 100 436 124
421 105 429 121
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
412 54 431 78
417 59 425 75
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
226 329 245 353
231 335 239 351
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
178 339 205 363
183 345 199 361
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
179 287 200 311
185 293 193 309
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
100 56 121 80
106 62 114 78
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
100 103 123 127
107 108 115 124
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
150 95 173 119
157 100 165 116
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
186 86 233 110
193 91 225 107
4 Y=A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
94 160 115 184
100 166 108 182
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
94 210 117 234
101 215 109 231
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
138 199 161 223
145 204 153 220
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
178 172 197 216
183 177 191 209
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
182 217 201 261
187 223 195 255
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
229 205 250 249
235 211 243 243
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
275 210 322 234
282 215 314 231
4 Y=AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
78 259 99 283
84 265 92 281
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
78 307 101 331
85 312 93 328
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
124 296 147 320
131 301 139 317
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
78 334 97 378
83 339 91 371
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
75 385 96 429
81 390 89 422
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
128 376 147 400
133 381 141 397
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
131 169 186 213
138 175 178 207
5 (AB)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
264 328 319 352
271 334 311 350
5 Y=A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
124 268 155 292
131 273 147 289
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
127 343 158 367
134 349 150 365
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
512 85 559 109
519 90 551 106
4 Y=A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
466 203 497 227
473 209 489 225
2 B'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
467 128 498 152
474 133 490 149
2 A'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
619 188 666 212
626 193 658 209
4 Y=AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
608 331 663 355
615 337 655 353
5 Y=A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
460 296 523 320
467 302 515 318
6 (A+B)'
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
