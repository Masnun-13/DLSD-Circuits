CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 40 1 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
41 D:\LEKHAPORA\FUBAR\Circuit Killer\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 78 96 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 L1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9466 0 0
2
44114.9 2
0
13 Logic Switch~
5 109 250 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 CLR1
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3266 0 0
2
44114.9 1
0
13 Logic Switch~
5 107 128 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 PRE1
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7693 0 0
2
44114.9 0
0
13 Logic Switch~
5 44 528 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 M
-2 -26 5 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3723 0 0
2
44114.9 12
0
13 Logic Switch~
5 78 627 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 L9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
44114.9 11
0
13 Logic Switch~
5 109 781 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 CLR3
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6263 0 0
2
44114.9 10
0
13 Logic Switch~
5 107 659 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 PRE3
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4900 0 0
2
44114.9 9
0
13 Logic Switch~
5 58 347 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 L8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8783 0 0
2
44114.9 6
0
13 Logic Switch~
5 89 498 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 CLR2
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3221 0 0
2
44114.9 5
0
13 Logic Switch~
5 123 376 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
4 PRE2
-12 -27 16 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3215 0 0
2
44114.9 4
0
7 Pulser~
4 76 174 0 10 12
0 28 2 29 2 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7903 0 0
2
44114.9 9
0
14 Logic Display~
6 273 73 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7121 0 0
2
44114.9 8
0
14 Logic Display~
6 488 71 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
44114.9 7
0
14 Logic Display~
6 709 68 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
44114.9 6
0
5 4027~
219 212 192 0 7 32
0 3 8 2 8 4 30 7
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
7804 0 0
2
44114.9 5
0
5 4027~
219 423 192 0 7 32
0 3 8 7 8 4 31 6
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 9 0
1 U
5523 0 0
2
44114.9 4
0
5 4027~
219 617 192 0 7 32
0 3 8 6 8 4 32 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 9 0
1 U
3330 0 0
2
44114.9 3
0
9 2-In XOR~
219 525 695 0 3 22
0 12 11 9
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3465 0 0
2
44114.9 8
0
9 2-In XOR~
219 309 696 0 3 22
0 13 11 10
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
8396 0 0
2
44114.9 7
0
7 Pulser~
4 76 705 0 10 12
0 33 14 34 14 0 0 5 5 1
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3685 0 0
2
44114.9 6
0
14 Logic Display~
6 273 604 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
44114.9 5
0
14 Logic Display~
6 488 602 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
44114.9 4
0
14 Logic Display~
6 709 599 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
44114.9 3
0
5 4027~
219 212 723 0 7 32
0 15 18 14 18 16 35 13
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
9156 0 0
2
44114.9 2
0
5 4027~
219 423 723 0 7 32
0 15 18 10 18 16 36 12
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U4A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 8 0
1 U
5776 0 0
2
44114.9 1
0
5 4027~
219 617 723 0 7 32
0 15 18 9 18 16 37 17
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U6A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 10 0
1 U
7207 0 0
2
44114.9 0
0
14 Logic Display~
6 690 317 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
44114.9 22
0
14 Logic Display~
6 469 319 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
44114.9 21
0
7 Pulser~
4 56 425 0 10 12
0 27 38 27 39 0 0 5 5 1
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
754 0 0
2
44114.9 20
0
14 Logic Display~
6 283 314 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9767 0 0
2
44114.9 19
0
5 4027~
219 192 443 0 7 32
0 19 26 27 26 20 22 25
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U7B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 11 0
1 U
7978 0 0
2
44114.9 18
0
5 4027~
219 403 443 0 7 32
0 19 26 22 26 20 21 24
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U7A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 11 0
1 U
3142 0 0
2
44114.9 17
0
5 4027~
219 597 443 0 7 32
0 19 26 21 26 20 40 23
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U6B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 10 0
1 U
3284 0 0
2
44114.9 16
0
61
0 4 2 0 0 8208 0 0 11 2 0 3
120 165
120 174
106 174
2 3 2 0 0 12432 0 11 15 0 0 6
46 174
37 174
37 141
120 141
120 165
188 165
0 1 3 0 0 4112 0 0 17 4 0 3
423 128
617 128
617 135
0 1 3 0 0 4240 0 0 16 5 0 3
212 128
423 128
423 135
1 1 3 0 0 16 0 3 15 0 0 3
119 128
212 128
212 135
0 5 4 0 0 4112 0 0 17 7 0 3
423 250
617 250
617 198
0 5 4 0 0 4240 0 0 16 8 0 3
212 250
423 250
423 198
1 5 4 0 0 16 0 2 15 0 0 3
121 250
212 250
212 198
7 1 5 0 0 8336 0 17 14 0 0 3
641 156
709 156
709 86
0 3 6 0 0 12304 0 0 17 11 0 4
487 156
530 156
530 165
593 165
7 1 6 0 0 8336 0 16 13 0 0 3
447 156
488 156
488 89
0 3 7 0 0 12432 0 0 16 13 0 4
272 156
334 156
334 165
399 165
7 1 7 0 0 16 0 15 12 0 0 3
236 156
273 156
273 91
0 4 8 0 0 4112 0 0 17 15 0 3
578 156
578 174
593 174
0 2 8 0 0 4112 0 0 17 17 0 4
389 96
578 96
578 156
593 156
0 4 8 0 0 16 0 0 16 17 0 3
390 156
390 174
399 174
0 2 8 0 0 4240 0 0 16 19 0 4
178 96
390 96
390 156
399 156
0 4 8 0 0 16 0 0 15 19 0 3
179 155
179 174
188 174
1 2 8 0 0 16 0 1 15 0 0 4
90 96
179 96
179 156
188 156
3 3 9 0 0 8320 0 18 26 0 0 3
558 695
558 696
593 696
3 3 10 0 0 4224 0 25 19 0 0 2
399 696
342 696
0 2 11 0 0 8320 0 0 18 23 0 5
271 705
271 748
480 748
480 704
509 704
1 2 11 0 0 0 0 4 19 0 0 4
56 528
255 528
255 705
293 705
0 1 12 0 0 8192 0 0 18 35 0 3
488 687
488 686
509 686
0 1 13 0 0 4096 0 0 19 36 0 2
273 687
293 687
0 4 14 0 0 8192 0 0 20 27 0 3
120 696
120 705
106 705
2 3 14 0 0 12416 0 20 24 0 0 6
46 705
37 705
37 672
120 672
120 696
188 696
0 1 15 0 0 4096 0 0 26 29 0 3
423 659
617 659
617 666
0 1 15 0 0 4224 0 0 25 30 0 3
212 659
423 659
423 666
1 1 15 0 0 0 0 7 24 0 0 3
119 659
212 659
212 666
0 5 16 0 0 4096 0 0 26 32 0 3
423 781
617 781
617 729
0 5 16 0 0 4224 0 0 25 33 0 3
212 781
423 781
423 729
1 5 16 0 0 0 0 6 24 0 0 3
121 781
212 781
212 729
7 1 17 0 0 8320 0 26 23 0 0 3
641 687
709 687
709 617
7 1 12 0 0 8320 0 25 22 0 0 3
447 687
488 687
488 620
7 1 13 0 0 8320 0 24 21 0 0 3
236 687
273 687
273 622
0 4 18 0 0 4096 0 0 26 38 0 3
578 687
578 705
593 705
0 2 18 0 0 4096 0 0 26 40 0 4
389 627
578 627
578 687
593 687
0 4 18 0 0 0 0 0 25 40 0 3
390 687
390 705
399 705
0 2 18 0 0 4224 0 0 25 42 0 4
178 627
390 627
390 687
399 687
0 4 18 0 0 0 0 0 24 42 0 3
179 686
179 705
188 705
1 2 18 0 0 0 0 5 24 0 0 4
90 627
179 627
179 687
188 687
0 1 19 0 0 8192 0 0 31 45 0 3
191 376
192 376
192 386
0 1 19 0 0 0 0 0 32 45 0 2
403 376
403 386
1 1 19 0 0 4224 0 10 33 0 0 3
135 376
597 376
597 386
0 5 20 0 0 4096 0 0 33 47 0 3
403 498
597 498
597 449
0 5 20 0 0 4224 0 0 32 48 0 3
192 498
403 498
403 449
1 5 20 0 0 0 0 9 31 0 0 3
101 498
192 498
192 449
6 3 21 0 0 4224 0 32 33 0 0 4
433 425
539 425
539 416
573 416
6 3 22 0 0 4224 0 31 32 0 0 4
222 425
329 425
329 416
379 416
7 1 23 0 0 8320 0 33 27 0 0 3
621 407
690 407
690 335
7 1 24 0 0 8320 0 32 28 0 0 3
427 407
469 407
469 337
7 1 25 0 0 8320 0 31 30 0 0 3
216 407
283 407
283 332
0 4 26 0 0 4096 0 0 33 55 0 3
558 407
558 425
573 425
0 2 26 0 0 4096 0 0 33 57 0 4
369 347
558 347
558 407
573 407
0 4 26 0 0 0 0 0 32 57 0 3
370 407
370 425
379 425
0 2 26 0 0 4224 0 0 32 59 0 4
158 347
370 347
370 407
379 407
0 4 26 0 0 0 0 0 31 59 0 3
159 406
159 425
168 425
1 2 26 0 0 0 0 8 31 0 0 4
70 347
159 347
159 407
168 407
1 0 27 0 0 12288 0 29 0 0 61 5
32 416
23 416
23 390
94 390
94 416
3 3 27 0 0 4224 0 29 31 0 0 2
80 416
168 416
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
